module AXI_FULL_MASTER(

);




endmodule
