module ysyx_20020207_CSRU(
  input clock, wen, decode_valid, ctrl_valid,
  input[2:0] csr_ctrl,
  input [11:0]csr_addr,
  input[31:0] wdata, pc,
  input lsu_ready,
  output reg[31:0] rdata, upc
);
`define MRET 3'b001
`define ECALL 3'b010
`define EBREAK 3'b011
`define CSRW 3'b100
  localparam MSTATUS = 2'b00;
  localparam MTVEC = 2'b01;
  localparam MEPC = 2'b10;
  localparam MCAUSE = 2'b11;
  reg[31:0] csr [3:0];
  reg[11:0] addr;
  always@(posedge clock)begin
    if(decode_valid) addr <= csr_addr;
  end
  
  reg[2:0] ctrl;
  always@(posedge clock)begin
    if(ctrl_valid) ctrl <= csr_ctrl;
  end

  reg[1:0] addr_map;
  always@(*)begin
    case(addr)
      12'h300: begin addr_map = MSTATUS; end
      12'h305: begin addr_map = MTVEC; end
      12'h341: begin addr_map = MEPC; end
      12'h342: begin addr_map = MCAUSE; end
      default: begin addr_map = 2'b00; end
    endcase
  end

   always @(posedge clock) begin
     if (lsu_ready && wen) begin
      case(ctrl)
        `CSRW:  begin csr[addr_map] <= wdata; end
        `ECALL: begin csr[MEPC] <= pc; csr[MCAUSE] <= 32'h0b; end
        default: begin end
      endcase
    end
  end

  always@(*)begin
    case(ctrl)
      `MRET:  begin upc = csr[MEPC]; end
      `ECALL: begin upc = csr[MTVEC]; end
      default begin upc = 0; end
    endcase
    if(addr_map == MSTATUS) rdata = 32'h1800;
    else rdata = csr[addr_map];
  end
  endmodule
