//Generate the verilog at 2024-05-05T20:53:09
module top (
clk,
exit,
jump,
lsu_finish,
mem_wen,
read_valid,
rst,
inst,
pc,
result,
upc
);

input clk ;
output exit ;
output jump ;
output lsu_finish ;
output mem_wen ;
input read_valid ;
input rst ;
output [31:0] inst ;
output [31:0] pc ;
output [31:0] result ;
output [31:0] upc ;

wire _000_ ;
wire _001_ ;
wire _002_ ;
wire _003_ ;
wire _004_ ;
wire _005_ ;
wire _006_ ;
wire _007_ ;
wire _008_ ;
wire _009_ ;
wire _010_ ;
wire _011_ ;
wire _012_ ;
wire _013_ ;
wire _014_ ;
wire _015_ ;
wire _016_ ;
wire _017_ ;
wire _018_ ;
wire _019_ ;
wire _020_ ;
wire _021_ ;
wire _022_ ;
wire _023_ ;
wire _024_ ;
wire _025_ ;
wire _026_ ;
wire _027_ ;
wire _028_ ;
wire _029_ ;
wire _030_ ;
wire _031_ ;
wire _032_ ;
wire _033_ ;
wire _034_ ;
wire _035_ ;
wire _036_ ;
wire _037_ ;
wire _038_ ;
wire _039_ ;
wire _040_ ;
wire _041_ ;
wire _042_ ;
wire _043_ ;
wire _044_ ;
wire _045_ ;
wire _046_ ;
wire _047_ ;
wire _048_ ;
wire _049_ ;
wire _050_ ;
wire _051_ ;
wire _052_ ;
wire _053_ ;
wire _054_ ;
wire _055_ ;
wire _056_ ;
wire _057_ ;
wire _058_ ;
wire _059_ ;
wire _060_ ;
wire _061_ ;
wire _062_ ;
wire _063_ ;
wire _064_ ;
wire _065_ ;
wire _066_ ;
wire _067_ ;
wire _068_ ;
wire _069_ ;
wire _070_ ;
wire _071_ ;
wire _072_ ;
wire _073_ ;
wire _074_ ;
wire _075_ ;
wire _076_ ;
wire _077_ ;
wire _078_ ;
wire _079_ ;
wire _080_ ;
wire _081_ ;
wire _082_ ;
wire _083_ ;
wire _084_ ;
wire _085_ ;
wire _086_ ;
wire _087_ ;
wire _088_ ;
wire _089_ ;
wire _090_ ;
wire _091_ ;
wire _092_ ;
wire _093_ ;
wire _094_ ;
wire _095_ ;
wire _096_ ;
wire _097_ ;
wire _098_ ;
wire _099_ ;
wire _100_ ;
wire _101_ ;
wire _102_ ;
wire _103_ ;
wire _104_ ;
wire _105_ ;
wire _106_ ;
wire _107_ ;
wire _108_ ;
wire _109_ ;
wire _110_ ;
wire _111_ ;
wire _112_ ;
wire _113_ ;
wire _114_ ;
wire _115_ ;
wire _116_ ;
wire _117_ ;
wire _118_ ;
wire _119_ ;
wire _120_ ;
wire _121_ ;
wire _122_ ;
wire _123_ ;
wire _124_ ;
wire _125_ ;
wire _126_ ;
wire _127_ ;
wire _128_ ;
wire _129_ ;
wire _130_ ;
wire _131_ ;
wire _132_ ;
wire _133_ ;
wire _134_ ;
wire _135_ ;
wire _136_ ;
wire _137_ ;
wire _138_ ;
wire _139_ ;
wire _140_ ;
wire _141_ ;
wire _142_ ;
wire _143_ ;
wire _144_ ;
wire _145_ ;
wire _146_ ;
wire _147_ ;
wire _148_ ;
wire _149_ ;
wire _150_ ;
wire _151_ ;
wire _152_ ;
wire _153_ ;
wire _154_ ;
wire _155_ ;
wire _156_ ;
wire _157_ ;
wire _158_ ;
wire _159_ ;
wire _160_ ;
wire _161_ ;
wire _162_ ;
wire _163_ ;
wire _164_ ;
wire _165_ ;
wire _166_ ;
wire _167_ ;
wire _168_ ;
wire _169_ ;
wire _170_ ;
wire _171_ ;
wire _172_ ;
wire _173_ ;
wire _174_ ;
wire _175_ ;
wire _176_ ;
wire _177_ ;
wire _178_ ;
wire _179_ ;
wire _180_ ;
wire _181_ ;
wire _182_ ;
wire _183_ ;
wire _184_ ;
wire _185_ ;
wire _186_ ;
wire _187_ ;
wire _188_ ;
wire _189_ ;
wire _190_ ;
wire _191_ ;
wire _192_ ;
wire _193_ ;
wire _194_ ;
wire _195_ ;
wire _196_ ;
wire _197_ ;
wire _198_ ;
wire _199_ ;
wire _200_ ;
wire _201_ ;
wire _202_ ;
wire _203_ ;
wire _204_ ;
wire _205_ ;
wire _206_ ;
wire _207_ ;
wire _208_ ;
wire _209_ ;
wire _210_ ;
wire _211_ ;
wire _212_ ;
wire _213_ ;
wire _214_ ;
wire _215_ ;
wire _216_ ;
wire _217_ ;
wire _218_ ;
wire _219_ ;
wire _220_ ;
wire _221_ ;
wire _222_ ;
wire _223_ ;
wire _224_ ;
wire _225_ ;
wire _226_ ;
wire _227_ ;
wire _228_ ;
wire _229_ ;
wire _230_ ;
wire _231_ ;
wire _232_ ;
wire _233_ ;
wire _234_ ;
wire _235_ ;
wire _236_ ;
wire _237_ ;
wire _238_ ;
wire _239_ ;
wire _240_ ;
wire _241_ ;
wire _242_ ;
wire _243_ ;
wire _244_ ;
wire _245_ ;
wire _246_ ;
wire _247_ ;
wire _248_ ;
wire _249_ ;
wire _250_ ;
wire _251_ ;
wire _252_ ;
wire _253_ ;
wire _254_ ;
wire _255_ ;
wire _256_ ;
wire _257_ ;
wire _258_ ;
wire _259_ ;
wire _260_ ;
wire _261_ ;
wire _262_ ;
wire _263_ ;
wire _264_ ;
wire _265_ ;
wire _266_ ;
wire _267_ ;
wire _268_ ;
wire _269_ ;
wire _270_ ;
wire _271_ ;
wire _272_ ;
wire _273_ ;
wire _274_ ;
wire _275_ ;
wire _276_ ;
wire _277_ ;
wire _278_ ;
wire _279_ ;
wire _280_ ;
wire _281_ ;
wire _282_ ;
wire _283_ ;
wire _284_ ;
wire _285_ ;
wire _286_ ;
wire _287_ ;
wire _288_ ;
wire _289_ ;
wire _290_ ;
wire _291_ ;
wire _292_ ;
wire _293_ ;
wire _294_ ;
wire _295_ ;
wire _296_ ;
wire _297_ ;
wire _298_ ;
wire _299_ ;
wire _300_ ;
wire _301_ ;
wire _302_ ;
wire _303_ ;
wire _304_ ;
wire _305_ ;
wire _306_ ;
wire _307_ ;
wire _308_ ;
wire _309_ ;
wire _310_ ;
wire _311_ ;
wire _312_ ;
wire _313_ ;
wire _314_ ;
wire _315_ ;
wire _316_ ;
wire _317_ ;
wire _318_ ;
wire _319_ ;
wire _320_ ;
wire _321_ ;
wire _322_ ;
wire _323_ ;
wire _324_ ;
wire _325_ ;
wire _326_ ;
wire _327_ ;
wire _328_ ;
wire _329_ ;
wire _330_ ;
wire _331_ ;
wire _332_ ;
wire _333_ ;
wire _334_ ;
wire _335_ ;
wire _336_ ;
wire _337_ ;
wire _338_ ;
wire _339_ ;
wire _340_ ;
wire _341_ ;
wire _342_ ;
wire _343_ ;
wire _344_ ;
wire _345_ ;
wire _346_ ;
wire _347_ ;
wire _348_ ;
wire _349_ ;
wire _350_ ;
wire _351_ ;
wire CF ;
wire OF ;
wire ZF ;
wire \alu_a[0] ;
wire \alu_a[10] ;
wire \alu_a[11] ;
wire \alu_a[12] ;
wire \alu_a[13] ;
wire \alu_a[14] ;
wire \alu_a[15] ;
wire \alu_a[16] ;
wire \alu_a[17] ;
wire \alu_a[18] ;
wire \alu_a[19] ;
wire \alu_a[1] ;
wire \alu_a[20] ;
wire \alu_a[21] ;
wire \alu_a[22] ;
wire \alu_a[23] ;
wire \alu_a[24] ;
wire \alu_a[25] ;
wire \alu_a[26] ;
wire \alu_a[27] ;
wire \alu_a[28] ;
wire \alu_a[29] ;
wire \alu_a[2] ;
wire \alu_a[30] ;
wire \alu_a[31] ;
wire \alu_a[3] ;
wire \alu_a[4] ;
wire \alu_a[5] ;
wire \alu_a[6] ;
wire \alu_a[7] ;
wire \alu_a[8] ;
wire \alu_a[9] ;
wire \alu_b[0] ;
wire \alu_b[10] ;
wire \alu_b[11] ;
wire \alu_b[12] ;
wire \alu_b[13] ;
wire \alu_b[14] ;
wire \alu_b[15] ;
wire \alu_b[16] ;
wire \alu_b[17] ;
wire \alu_b[18] ;
wire \alu_b[19] ;
wire \alu_b[1] ;
wire \alu_b[20] ;
wire \alu_b[21] ;
wire \alu_b[22] ;
wire \alu_b[23] ;
wire \alu_b[24] ;
wire \alu_b[25] ;
wire \alu_b[26] ;
wire \alu_b[27] ;
wire \alu_b[28] ;
wire \alu_b[29] ;
wire \alu_b[2] ;
wire \alu_b[30] ;
wire \alu_b[31] ;
wire \alu_b[3] ;
wire \alu_b[4] ;
wire \alu_b[5] ;
wire \alu_b[6] ;
wire \alu_b[7] ;
wire \alu_b[8] ;
wire \alu_b[9] ;
wire \alu_ctl[0] ;
wire \alu_ctl[1] ;
wire \alu_ctl[2] ;
wire \alu_ctl[3] ;
wire \alu_result[0] ;
wire \alu_result[10] ;
wire \alu_result[11] ;
wire \alu_result[12] ;
wire \alu_result[13] ;
wire \alu_result[14] ;
wire \alu_result[15] ;
wire \alu_result[16] ;
wire \alu_result[17] ;
wire \alu_result[18] ;
wire \alu_result[19] ;
wire \alu_result[1] ;
wire \alu_result[20] ;
wire \alu_result[21] ;
wire \alu_result[22] ;
wire \alu_result[23] ;
wire \alu_result[24] ;
wire \alu_result[25] ;
wire \alu_result[26] ;
wire \alu_result[27] ;
wire \alu_result[28] ;
wire \alu_result[29] ;
wire \alu_result[2] ;
wire \alu_result[30] ;
wire \alu_result[31] ;
wire \alu_result[3] ;
wire \alu_result[4] ;
wire \alu_result[5] ;
wire \alu_result[6] ;
wire \alu_result[7] ;
wire \alu_result[8] ;
wire \alu_result[9] ;
wire alu_sign ;
wire alu_sub ;
wire \araddr[0] ;
wire \araddr[10] ;
wire \araddr[11] ;
wire \araddr[12] ;
wire \araddr[13] ;
wire \araddr[14] ;
wire \araddr[15] ;
wire \araddr[16] ;
wire \araddr[17] ;
wire \araddr[18] ;
wire \araddr[19] ;
wire \araddr[1] ;
wire \araddr[20] ;
wire \araddr[21] ;
wire \araddr[22] ;
wire \araddr[23] ;
wire \araddr[24] ;
wire \araddr[25] ;
wire \araddr[26] ;
wire \araddr[27] ;
wire \araddr[28] ;
wire \araddr[29] ;
wire \araddr[2] ;
wire \araddr[30] ;
wire \araddr[31] ;
wire \araddr[3] ;
wire \araddr[4] ;
wire \araddr[5] ;
wire \araddr[6] ;
wire \araddr[7] ;
wire \araddr[8] ;
wire \araddr[9] ;
wire arready ;
wire arvalid ;
wire \awaddr[0] ;
wire \awaddr[10] ;
wire \awaddr[11] ;
wire \awaddr[12] ;
wire \awaddr[13] ;
wire \awaddr[14] ;
wire \awaddr[15] ;
wire \awaddr[16] ;
wire \awaddr[17] ;
wire \awaddr[18] ;
wire \awaddr[19] ;
wire \awaddr[1] ;
wire \awaddr[20] ;
wire \awaddr[21] ;
wire \awaddr[22] ;
wire \awaddr[23] ;
wire \awaddr[24] ;
wire \awaddr[25] ;
wire \awaddr[26] ;
wire \awaddr[27] ;
wire \awaddr[28] ;
wire \awaddr[29] ;
wire \awaddr[2] ;
wire \awaddr[30] ;
wire \awaddr[31] ;
wire \awaddr[3] ;
wire \awaddr[4] ;
wire \awaddr[5] ;
wire \awaddr[6] ;
wire \awaddr[7] ;
wire \awaddr[8] ;
wire \awaddr[9] ;
wire awready ;
wire awvalid ;
wire branch ;
wire bready ;
wire \bresp[0] ;
wire \bresp[1] ;
wire bvalid ;
wire clk ;
wire \csr_ctl[0] ;
wire \csr_ctl[1] ;
wire \csr_ctl[2] ;
wire \csr_rdata[0] ;
wire \csr_rdata[10] ;
wire \csr_rdata[11] ;
wire \csr_rdata[12] ;
wire \csr_rdata[13] ;
wire \csr_rdata[14] ;
wire \csr_rdata[15] ;
wire \csr_rdata[16] ;
wire \csr_rdata[17] ;
wire \csr_rdata[18] ;
wire \csr_rdata[19] ;
wire \csr_rdata[1] ;
wire \csr_rdata[20] ;
wire \csr_rdata[21] ;
wire \csr_rdata[22] ;
wire \csr_rdata[23] ;
wire \csr_rdata[24] ;
wire \csr_rdata[25] ;
wire \csr_rdata[26] ;
wire \csr_rdata[27] ;
wire \csr_rdata[28] ;
wire \csr_rdata[29] ;
wire \csr_rdata[2] ;
wire \csr_rdata[30] ;
wire \csr_rdata[31] ;
wire \csr_rdata[3] ;
wire \csr_rdata[4] ;
wire \csr_rdata[5] ;
wire \csr_rdata[6] ;
wire \csr_rdata[7] ;
wire \csr_rdata[8] ;
wire \csr_rdata[9] ;
wire \csr_upc[0] ;
wire \csr_upc[10] ;
wire \csr_upc[11] ;
wire \csr_upc[12] ;
wire \csr_upc[13] ;
wire \csr_upc[14] ;
wire \csr_upc[15] ;
wire \csr_upc[16] ;
wire \csr_upc[17] ;
wire \csr_upc[18] ;
wire \csr_upc[19] ;
wire \csr_upc[1] ;
wire \csr_upc[20] ;
wire \csr_upc[21] ;
wire \csr_upc[22] ;
wire \csr_upc[23] ;
wire \csr_upc[24] ;
wire \csr_upc[25] ;
wire \csr_upc[26] ;
wire \csr_upc[27] ;
wire \csr_upc[28] ;
wire \csr_upc[29] ;
wire \csr_upc[2] ;
wire \csr_upc[30] ;
wire \csr_upc[31] ;
wire \csr_upc[3] ;
wire \csr_upc[4] ;
wire \csr_upc[5] ;
wire \csr_upc[6] ;
wire \csr_upc[7] ;
wire \csr_upc[8] ;
wire \csr_upc[9] ;
wire csr_wen ;
wire exit ;
wire exu_jump ;
wire \exu_upc[0] ;
wire \exu_upc[10] ;
wire \exu_upc[11] ;
wire \exu_upc[12] ;
wire \exu_upc[13] ;
wire \exu_upc[14] ;
wire \exu_upc[15] ;
wire \exu_upc[16] ;
wire \exu_upc[17] ;
wire \exu_upc[18] ;
wire \exu_upc[19] ;
wire \exu_upc[1] ;
wire \exu_upc[20] ;
wire \exu_upc[21] ;
wire \exu_upc[22] ;
wire \exu_upc[23] ;
wire \exu_upc[24] ;
wire \exu_upc[25] ;
wire \exu_upc[26] ;
wire \exu_upc[27] ;
wire \exu_upc[28] ;
wire \exu_upc[29] ;
wire \exu_upc[2] ;
wire \exu_upc[30] ;
wire \exu_upc[31] ;
wire \exu_upc[3] ;
wire \exu_upc[4] ;
wire \exu_upc[5] ;
wire \exu_upc[6] ;
wire \exu_upc[7] ;
wire \exu_upc[8] ;
wire \exu_upc[9] ;
wire \func[0] ;
wire \func[1] ;
wire \func[2] ;
wire \ifu_araddr[0] ;
wire \ifu_araddr[10] ;
wire \ifu_araddr[11] ;
wire \ifu_araddr[12] ;
wire \ifu_araddr[13] ;
wire \ifu_araddr[14] ;
wire \ifu_araddr[15] ;
wire \ifu_araddr[16] ;
wire \ifu_araddr[17] ;
wire \ifu_araddr[18] ;
wire \ifu_araddr[19] ;
wire \ifu_araddr[1] ;
wire \ifu_araddr[20] ;
wire \ifu_araddr[21] ;
wire \ifu_araddr[22] ;
wire \ifu_araddr[23] ;
wire \ifu_araddr[24] ;
wire \ifu_araddr[25] ;
wire \ifu_araddr[26] ;
wire \ifu_araddr[27] ;
wire \ifu_araddr[28] ;
wire \ifu_araddr[29] ;
wire \ifu_araddr[2] ;
wire \ifu_araddr[30] ;
wire \ifu_araddr[31] ;
wire \ifu_araddr[3] ;
wire \ifu_araddr[4] ;
wire \ifu_araddr[5] ;
wire \ifu_araddr[6] ;
wire \ifu_araddr[7] ;
wire \ifu_araddr[8] ;
wire \ifu_araddr[9] ;
wire ifu_arready ;
wire ifu_arvalid ;
wire ifu_awready ;
wire \ifu_bresp[0] ;
wire \ifu_bresp[1] ;
wire ifu_bvalid ;
wire \ifu_rdata[0] ;
wire \ifu_rdata[10] ;
wire \ifu_rdata[11] ;
wire \ifu_rdata[12] ;
wire \ifu_rdata[13] ;
wire \ifu_rdata[14] ;
wire \ifu_rdata[15] ;
wire \ifu_rdata[16] ;
wire \ifu_rdata[17] ;
wire \ifu_rdata[18] ;
wire \ifu_rdata[19] ;
wire \ifu_rdata[1] ;
wire \ifu_rdata[20] ;
wire \ifu_rdata[21] ;
wire \ifu_rdata[22] ;
wire \ifu_rdata[23] ;
wire \ifu_rdata[24] ;
wire \ifu_rdata[25] ;
wire \ifu_rdata[26] ;
wire \ifu_rdata[27] ;
wire \ifu_rdata[28] ;
wire \ifu_rdata[29] ;
wire \ifu_rdata[2] ;
wire \ifu_rdata[30] ;
wire \ifu_rdata[31] ;
wire \ifu_rdata[3] ;
wire \ifu_rdata[4] ;
wire \ifu_rdata[5] ;
wire \ifu_rdata[6] ;
wire \ifu_rdata[7] ;
wire \ifu_rdata[8] ;
wire \ifu_rdata[9] ;
wire ifu_rready ;
wire \ifu_rresp[0] ;
wire \ifu_rresp[1] ;
wire ifu_rvalid ;
wire ifu_wready ;
wire \imm[0] ;
wire \imm[10] ;
wire \imm[11] ;
wire \imm[12] ;
wire \imm[13] ;
wire \imm[14] ;
wire \imm[15] ;
wire \imm[16] ;
wire \imm[17] ;
wire \imm[18] ;
wire \imm[19] ;
wire \imm[1] ;
wire \imm[20] ;
wire \imm[21] ;
wire \imm[22] ;
wire \imm[23] ;
wire \imm[24] ;
wire \imm[25] ;
wire \imm[26] ;
wire \imm[27] ;
wire \imm[28] ;
wire \imm[29] ;
wire \imm[2] ;
wire \imm[30] ;
wire \imm[31] ;
wire \imm[3] ;
wire \imm[4] ;
wire \imm[5] ;
wire \imm[6] ;
wire \imm[7] ;
wire \imm[8] ;
wire \imm[9] ;
wire \inst[0] ;
wire \inst[1] ;
wire \inst[2] ;
wire \inst[3] ;
wire \inst[4] ;
wire \inst[5] ;
wire \inst[6] ;
wire \inst[7] ;
wire \inst[8] ;
wire \inst[9] ;
wire \inst[10] ;
wire \inst[11] ;
wire \inst[12] ;
wire \inst[13] ;
wire \inst[14] ;
wire \inst[15] ;
wire \inst[16] ;
wire \inst[17] ;
wire \inst[18] ;
wire \inst[19] ;
wire \inst[20] ;
wire \inst[21] ;
wire \inst[22] ;
wire \inst[23] ;
wire \inst[24] ;
wire \inst[25] ;
wire \inst[26] ;
wire \inst[27] ;
wire \inst[28] ;
wire \inst[29] ;
wire \inst[30] ;
wire \inst[31] ;
wire inst_valid ;
wire jump ;
wire \load_ctl[0] ;
wire \load_ctl[1] ;
wire \load_ctl[2] ;
wire \lsu_araddr[0] ;
wire \lsu_araddr[10] ;
wire \lsu_araddr[11] ;
wire \lsu_araddr[12] ;
wire \lsu_araddr[13] ;
wire \lsu_araddr[14] ;
wire \lsu_araddr[15] ;
wire \lsu_araddr[16] ;
wire \lsu_araddr[17] ;
wire \lsu_araddr[18] ;
wire \lsu_araddr[19] ;
wire \lsu_araddr[1] ;
wire \lsu_araddr[20] ;
wire \lsu_araddr[21] ;
wire \lsu_araddr[22] ;
wire \lsu_araddr[23] ;
wire \lsu_araddr[24] ;
wire \lsu_araddr[25] ;
wire \lsu_araddr[26] ;
wire \lsu_araddr[27] ;
wire \lsu_araddr[28] ;
wire \lsu_araddr[29] ;
wire \lsu_araddr[2] ;
wire \lsu_araddr[30] ;
wire \lsu_araddr[31] ;
wire \lsu_araddr[3] ;
wire \lsu_araddr[4] ;
wire \lsu_araddr[5] ;
wire \lsu_araddr[6] ;
wire \lsu_araddr[7] ;
wire \lsu_araddr[8] ;
wire \lsu_araddr[9] ;
wire lsu_arready ;
wire lsu_arvalid ;
wire \lsu_awaddr[0] ;
wire \lsu_awaddr[10] ;
wire \lsu_awaddr[11] ;
wire \lsu_awaddr[12] ;
wire \lsu_awaddr[13] ;
wire \lsu_awaddr[14] ;
wire \lsu_awaddr[15] ;
wire \lsu_awaddr[16] ;
wire \lsu_awaddr[17] ;
wire \lsu_awaddr[18] ;
wire \lsu_awaddr[19] ;
wire \lsu_awaddr[1] ;
wire \lsu_awaddr[20] ;
wire \lsu_awaddr[21] ;
wire \lsu_awaddr[22] ;
wire \lsu_awaddr[23] ;
wire \lsu_awaddr[24] ;
wire \lsu_awaddr[25] ;
wire \lsu_awaddr[26] ;
wire \lsu_awaddr[27] ;
wire \lsu_awaddr[28] ;
wire \lsu_awaddr[29] ;
wire \lsu_awaddr[2] ;
wire \lsu_awaddr[30] ;
wire \lsu_awaddr[31] ;
wire \lsu_awaddr[3] ;
wire \lsu_awaddr[4] ;
wire \lsu_awaddr[5] ;
wire \lsu_awaddr[6] ;
wire \lsu_awaddr[7] ;
wire \lsu_awaddr[8] ;
wire \lsu_awaddr[9] ;
wire lsu_awready ;
wire lsu_awvalid ;
wire lsu_bready ;
wire \lsu_bresp[0] ;
wire \lsu_bresp[1] ;
wire lsu_bvalid ;
wire lsu_finish ;
wire \lsu_rdata[0] ;
wire \lsu_rdata[10] ;
wire \lsu_rdata[11] ;
wire \lsu_rdata[12] ;
wire \lsu_rdata[13] ;
wire \lsu_rdata[14] ;
wire \lsu_rdata[15] ;
wire \lsu_rdata[16] ;
wire \lsu_rdata[17] ;
wire \lsu_rdata[18] ;
wire \lsu_rdata[19] ;
wire \lsu_rdata[1] ;
wire \lsu_rdata[20] ;
wire \lsu_rdata[21] ;
wire \lsu_rdata[22] ;
wire \lsu_rdata[23] ;
wire \lsu_rdata[24] ;
wire \lsu_rdata[25] ;
wire \lsu_rdata[26] ;
wire \lsu_rdata[27] ;
wire \lsu_rdata[28] ;
wire \lsu_rdata[29] ;
wire \lsu_rdata[2] ;
wire \lsu_rdata[30] ;
wire \lsu_rdata[31] ;
wire \lsu_rdata[3] ;
wire \lsu_rdata[4] ;
wire \lsu_rdata[5] ;
wire \lsu_rdata[6] ;
wire \lsu_rdata[7] ;
wire \lsu_rdata[8] ;
wire \lsu_rdata[9] ;
wire lsu_rready ;
wire \lsu_rresp[0] ;
wire \lsu_rresp[1] ;
wire lsu_rvalid ;
wire \lsu_wdata[0] ;
wire \lsu_wdata[10] ;
wire \lsu_wdata[11] ;
wire \lsu_wdata[12] ;
wire \lsu_wdata[13] ;
wire \lsu_wdata[14] ;
wire \lsu_wdata[15] ;
wire \lsu_wdata[16] ;
wire \lsu_wdata[17] ;
wire \lsu_wdata[18] ;
wire \lsu_wdata[19] ;
wire \lsu_wdata[1] ;
wire \lsu_wdata[20] ;
wire \lsu_wdata[21] ;
wire \lsu_wdata[22] ;
wire \lsu_wdata[23] ;
wire \lsu_wdata[24] ;
wire \lsu_wdata[25] ;
wire \lsu_wdata[26] ;
wire \lsu_wdata[27] ;
wire \lsu_wdata[28] ;
wire \lsu_wdata[29] ;
wire \lsu_wdata[2] ;
wire \lsu_wdata[30] ;
wire \lsu_wdata[31] ;
wire \lsu_wdata[3] ;
wire \lsu_wdata[4] ;
wire \lsu_wdata[5] ;
wire \lsu_wdata[6] ;
wire \lsu_wdata[7] ;
wire \lsu_wdata[8] ;
wire \lsu_wdata[9] ;
wire lsu_wready ;
wire \lsu_wstrb[0] ;
wire \lsu_wstrb[1] ;
wire \lsu_wstrb[2] ;
wire \lsu_wstrb[3] ;
wire \lsu_wstrb[4] ;
wire \lsu_wstrb[5] ;
wire \lsu_wstrb[6] ;
wire \lsu_wstrb[7] ;
wire lsu_wvalid ;
wire \mem_rdata[0] ;
wire \mem_rdata[10] ;
wire \mem_rdata[11] ;
wire \mem_rdata[12] ;
wire \mem_rdata[13] ;
wire \mem_rdata[14] ;
wire \mem_rdata[15] ;
wire \mem_rdata[16] ;
wire \mem_rdata[17] ;
wire \mem_rdata[18] ;
wire \mem_rdata[19] ;
wire \mem_rdata[1] ;
wire \mem_rdata[20] ;
wire \mem_rdata[21] ;
wire \mem_rdata[22] ;
wire \mem_rdata[23] ;
wire \mem_rdata[24] ;
wire \mem_rdata[25] ;
wire \mem_rdata[26] ;
wire \mem_rdata[27] ;
wire \mem_rdata[28] ;
wire \mem_rdata[29] ;
wire \mem_rdata[2] ;
wire \mem_rdata[30] ;
wire \mem_rdata[31] ;
wire \mem_rdata[3] ;
wire \mem_rdata[4] ;
wire \mem_rdata[5] ;
wire \mem_rdata[6] ;
wire \mem_rdata[7] ;
wire \mem_rdata[8] ;
wire \mem_rdata[9] ;
wire mem_ren ;
wire \mem_wdata[0] ;
wire \mem_wdata[10] ;
wire \mem_wdata[11] ;
wire \mem_wdata[12] ;
wire \mem_wdata[13] ;
wire \mem_wdata[14] ;
wire \mem_wdata[15] ;
wire \mem_wdata[16] ;
wire \mem_wdata[17] ;
wire \mem_wdata[18] ;
wire \mem_wdata[19] ;
wire \mem_wdata[1] ;
wire \mem_wdata[20] ;
wire \mem_wdata[21] ;
wire \mem_wdata[22] ;
wire \mem_wdata[23] ;
wire \mem_wdata[24] ;
wire \mem_wdata[25] ;
wire \mem_wdata[26] ;
wire \mem_wdata[27] ;
wire \mem_wdata[28] ;
wire \mem_wdata[29] ;
wire \mem_wdata[2] ;
wire \mem_wdata[30] ;
wire \mem_wdata[31] ;
wire \mem_wdata[3] ;
wire \mem_wdata[4] ;
wire \mem_wdata[5] ;
wire \mem_wdata[6] ;
wire \mem_wdata[7] ;
wire \mem_wdata[8] ;
wire \mem_wdata[9] ;
wire mem_wen ;
wire \op[0] ;
wire \op[1] ;
wire \op[2] ;
wire \op[3] ;
wire \op[4] ;
wire \op[5] ;
wire \op[6] ;
wire \pc[0] ;
wire \pc[1] ;
wire \pc[2] ;
wire \pc[3] ;
wire \pc[4] ;
wire \pc[5] ;
wire \pc[6] ;
wire \pc[7] ;
wire \pc[8] ;
wire \pc[9] ;
wire \pc[10] ;
wire \pc[11] ;
wire \pc[12] ;
wire \pc[13] ;
wire \pc[14] ;
wire \pc[15] ;
wire \pc[16] ;
wire \pc[17] ;
wire \pc[18] ;
wire \pc[19] ;
wire \pc[20] ;
wire \pc[21] ;
wire \pc[22] ;
wire \pc[23] ;
wire \pc[24] ;
wire \pc[25] ;
wire \pc[26] ;
wire \pc[27] ;
wire \pc[28] ;
wire \pc[29] ;
wire \pc[30] ;
wire \pc[31] ;
wire pc_wen ;
wire \rd[0] ;
wire \rd[1] ;
wire \rd[2] ;
wire \rd[3] ;
wire \rd[4] ;
wire \rdata[0] ;
wire \rdata[10] ;
wire \rdata[11] ;
wire \rdata[12] ;
wire \rdata[13] ;
wire \rdata[14] ;
wire \rdata[15] ;
wire \rdata[16] ;
wire \rdata[17] ;
wire \rdata[18] ;
wire \rdata[19] ;
wire \rdata[1] ;
wire \rdata[20] ;
wire \rdata[21] ;
wire \rdata[22] ;
wire \rdata[23] ;
wire \rdata[24] ;
wire \rdata[25] ;
wire \rdata[26] ;
wire \rdata[27] ;
wire \rdata[28] ;
wire \rdata[29] ;
wire \rdata[2] ;
wire \rdata[30] ;
wire \rdata[31] ;
wire \rdata[3] ;
wire \rdata[4] ;
wire \rdata[5] ;
wire \rdata[6] ;
wire \rdata[7] ;
wire \rdata[8] ;
wire \rdata[9] ;
wire read_valid ;
wire reg_wen ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;
wire \result[10] ;
wire \result[11] ;
wire \result[12] ;
wire \result[13] ;
wire \result[14] ;
wire \result[15] ;
wire \result[16] ;
wire \result[17] ;
wire \result[18] ;
wire \result[19] ;
wire \result[20] ;
wire \result[21] ;
wire \result[22] ;
wire \result[23] ;
wire \result[24] ;
wire \result[25] ;
wire \result[26] ;
wire \result[27] ;
wire \result[28] ;
wire \result[29] ;
wire \result[30] ;
wire \result[31] ;
wire \result_ctl[0] ;
wire \result_ctl[1] ;
wire rready ;
wire \rresp[0] ;
wire \rresp[1] ;
wire \rs1[0] ;
wire \rs1[1] ;
wire \rs1[2] ;
wire \rs1[3] ;
wire \rs1[4] ;
wire \rs2[0] ;
wire \rs2[1] ;
wire \rs2[2] ;
wire \rs2[3] ;
wire \rs2[4] ;
wire rst ;
wire rvalid ;
wire \src1[0] ;
wire \src1[10] ;
wire \src1[11] ;
wire \src1[12] ;
wire \src1[13] ;
wire \src1[14] ;
wire \src1[15] ;
wire \src1[16] ;
wire \src1[17] ;
wire \src1[18] ;
wire \src1[19] ;
wire \src1[1] ;
wire \src1[20] ;
wire \src1[21] ;
wire \src1[22] ;
wire \src1[23] ;
wire \src1[24] ;
wire \src1[25] ;
wire \src1[26] ;
wire \src1[27] ;
wire \src1[28] ;
wire \src1[29] ;
wire \src1[2] ;
wire \src1[30] ;
wire \src1[31] ;
wire \src1[3] ;
wire \src1[4] ;
wire \src1[5] ;
wire \src1[6] ;
wire \src1[7] ;
wire \src1[8] ;
wire \src1[9] ;
wire \upc[0] ;
wire \upc[1] ;
wire \upc[2] ;
wire \upc[3] ;
wire \upc[4] ;
wire \upc[5] ;
wire \upc[6] ;
wire \upc[7] ;
wire \upc[8] ;
wire \upc[9] ;
wire \upc[10] ;
wire \upc[11] ;
wire \upc[12] ;
wire \upc[13] ;
wire \upc[14] ;
wire \upc[15] ;
wire \upc[16] ;
wire \upc[17] ;
wire \upc[18] ;
wire \upc[19] ;
wire \upc[20] ;
wire \upc[21] ;
wire \upc[22] ;
wire \upc[23] ;
wire \upc[24] ;
wire \upc[25] ;
wire \upc[26] ;
wire \upc[27] ;
wire \upc[28] ;
wire \upc[29] ;
wire \upc[30] ;
wire \upc[31] ;
wire upc_ctl ;
wire \wdata[0] ;
wire \wdata[10] ;
wire \wdata[11] ;
wire \wdata[12] ;
wire \wdata[13] ;
wire \wdata[14] ;
wire \wdata[15] ;
wire \wdata[16] ;
wire \wdata[17] ;
wire \wdata[18] ;
wire \wdata[19] ;
wire \wdata[1] ;
wire \wdata[20] ;
wire \wdata[21] ;
wire \wdata[22] ;
wire \wdata[23] ;
wire \wdata[24] ;
wire \wdata[25] ;
wire \wdata[26] ;
wire \wdata[27] ;
wire \wdata[28] ;
wire \wdata[29] ;
wire \wdata[2] ;
wire \wdata[30] ;
wire \wdata[31] ;
wire \wdata[3] ;
wire \wdata[4] ;
wire \wdata[5] ;
wire \wdata[6] ;
wire \wdata[7] ;
wire \wdata[8] ;
wire \wdata[9] ;
wire \wmask[0] ;
wire \wmask[1] ;
wire \wmask[2] ;
wire \wmask[3] ;
wire \wmask[4] ;
wire \wmask[5] ;
wire \wmask[6] ;
wire \wmask[7] ;
wire wready ;
wire \wstrb[0] ;
wire \wstrb[1] ;
wire \wstrb[2] ;
wire \wstrb[3] ;
wire \wstrb[4] ;
wire \wstrb[5] ;
wire \wstrb[6] ;
wire \wstrb[7] ;
wire wvalid ;
wire \malu/_000_ ;
wire \malu/_001_ ;
wire \malu/_002_ ;
wire \malu/_003_ ;
wire \malu/_004_ ;
wire \malu/_005_ ;
wire \malu/_006_ ;
wire \malu/_007_ ;
wire \malu/_008_ ;
wire \malu/_009_ ;
wire \malu/_010_ ;
wire \malu/_011_ ;
wire \malu/_012_ ;
wire \malu/_013_ ;
wire \malu/_014_ ;
wire \malu/_015_ ;
wire \malu/_016_ ;
wire \malu/_017_ ;
wire \malu/_018_ ;
wire \malu/_019_ ;
wire \malu/_020_ ;
wire \malu/_021_ ;
wire \malu/_022_ ;
wire \malu/_023_ ;
wire \malu/_024_ ;
wire \malu/_025_ ;
wire \malu/_026_ ;
wire \malu/_027_ ;
wire \malu/_028_ ;
wire \malu/_029_ ;
wire \malu/_030_ ;
wire \malu/_031_ ;
wire \malu/_032_ ;
wire \malu/_033_ ;
wire \malu/_034_ ;
wire \malu/_035_ ;
wire \malu/_036_ ;
wire \malu/_037_ ;
wire \malu/_038_ ;
wire \malu/_039_ ;
wire \malu/_040_ ;
wire \malu/_041_ ;
wire \malu/_042_ ;
wire \malu/_043_ ;
wire \malu/_044_ ;
wire \malu/_045_ ;
wire \malu/_046_ ;
wire \malu/_047_ ;
wire \malu/_048_ ;
wire \malu/_049_ ;
wire \malu/_050_ ;
wire \malu/_051_ ;
wire \malu/_052_ ;
wire \malu/_053_ ;
wire \malu/_054_ ;
wire \malu/_055_ ;
wire \malu/_056_ ;
wire \malu/_057_ ;
wire \malu/_058_ ;
wire \malu/_059_ ;
wire \malu/_060_ ;
wire \malu/_061_ ;
wire \malu/_062_ ;
wire \malu/_063_ ;
wire \malu/_064_ ;
wire \malu/_065_ ;
wire \malu/_066_ ;
wire \malu/_067_ ;
wire \malu/_068_ ;
wire \malu/_069_ ;
wire \malu/_070_ ;
wire \malu/_071_ ;
wire \malu/_072_ ;
wire \malu/_073_ ;
wire \malu/_074_ ;
wire \malu/_075_ ;
wire \malu/_076_ ;
wire \malu/_077_ ;
wire \malu/_078_ ;
wire \malu/_079_ ;
wire \malu/_080_ ;
wire \malu/_081_ ;
wire \malu/_082_ ;
wire \malu/_083_ ;
wire \malu/_084_ ;
wire \malu/_085_ ;
wire \malu/_086_ ;
wire \malu/_087_ ;
wire \malu/_088_ ;
wire \malu/_089_ ;
wire \malu/_090_ ;
wire \malu/_091_ ;
wire \malu/_092_ ;
wire \malu/_093_ ;
wire \malu/_094_ ;
wire \malu/_095_ ;
wire \malu/_096_ ;
wire \malu/_097_ ;
wire \malu/_098_ ;
wire \malu/_099_ ;
wire \malu/_100_ ;
wire \malu/_101_ ;
wire \malu/_102_ ;
wire \malu/_103_ ;
wire \malu/_104_ ;
wire \malu/_105_ ;
wire \malu/_106_ ;
wire \malu/_107_ ;
wire \malu/_108_ ;
wire \malu/_109_ ;
wire \malu/_110_ ;
wire \malu/_111_ ;
wire \malu/_112_ ;
wire \malu/_113_ ;
wire \malu/_114_ ;
wire \malu/_115_ ;
wire \malu/_116_ ;
wire \malu/_117_ ;
wire \malu/_118_ ;
wire \malu/_119_ ;
wire \malu/_120_ ;
wire \malu/_121_ ;
wire \malu/_122_ ;
wire \malu/_123_ ;
wire \malu/_124_ ;
wire \malu/_125_ ;
wire \malu/_126_ ;
wire \malu/_127_ ;
wire \malu/_128_ ;
wire \malu/_129_ ;
wire \malu/_130_ ;
wire \malu/_131_ ;
wire \malu/_132_ ;
wire \malu/_133_ ;
wire \malu/_134_ ;
wire \malu/_135_ ;
wire \malu/_136_ ;
wire \malu/_137_ ;
wire \malu/_138_ ;
wire \malu/_139_ ;
wire \malu/_140_ ;
wire \malu/_141_ ;
wire \malu/_142_ ;
wire \malu/_143_ ;
wire \malu/_144_ ;
wire \malu/_145_ ;
wire \malu/_146_ ;
wire \malu/_147_ ;
wire \malu/_148_ ;
wire \malu/_149_ ;
wire \malu/_150_ ;
wire \malu/_151_ ;
wire \malu/_152_ ;
wire \malu/_153_ ;
wire \malu/_154_ ;
wire \malu/_155_ ;
wire \malu/_156_ ;
wire \malu/_157_ ;
wire \malu/_158_ ;
wire \malu/_159_ ;
wire \malu/_160_ ;
wire \malu/_161_ ;
wire \malu/_162_ ;
wire \malu/_163_ ;
wire \malu/_164_ ;
wire \malu/_165_ ;
wire \malu/_166_ ;
wire \malu/_167_ ;
wire \malu/_168_ ;
wire \malu/_169_ ;
wire \malu/_170_ ;
wire \malu/_171_ ;
wire \malu/_172_ ;
wire \malu/_173_ ;
wire \malu/_174_ ;
wire \malu/_175_ ;
wire \malu/_176_ ;
wire \malu/_177_ ;
wire \malu/_178_ ;
wire \malu/_179_ ;
wire \malu/_180_ ;
wire \malu/_181_ ;
wire \malu/_182_ ;
wire \malu/_183_ ;
wire \malu/_184_ ;
wire \malu/_185_ ;
wire \malu/_186_ ;
wire \malu/_187_ ;
wire \malu/_188_ ;
wire \malu/_189_ ;
wire \malu/_190_ ;
wire \malu/_191_ ;
wire \malu/_192_ ;
wire \malu/_193_ ;
wire \malu/_194_ ;
wire \malu/_195_ ;
wire \malu/_196_ ;
wire \malu/_197_ ;
wire \malu/_198_ ;
wire \malu/_199_ ;
wire \malu/_200_ ;
wire \malu/_201_ ;
wire \malu/_202_ ;
wire \malu/_203_ ;
wire \malu/_204_ ;
wire \malu/_205_ ;
wire \malu/_206_ ;
wire \malu/_207_ ;
wire \malu/_208_ ;
wire \malu/_209_ ;
wire \malu/_210_ ;
wire \malu/_211_ ;
wire \malu/_212_ ;
wire \malu/_213_ ;
wire \malu/_214_ ;
wire \malu/_215_ ;
wire \malu/_216_ ;
wire \malu/_217_ ;
wire \malu/_218_ ;
wire \malu/_219_ ;
wire \malu/_220_ ;
wire \malu/_221_ ;
wire \malu/_222_ ;
wire \malu/_223_ ;
wire \malu/_224_ ;
wire \malu/_225_ ;
wire \malu/_226_ ;
wire \malu/_227_ ;
wire \malu/_228_ ;
wire \malu/_229_ ;
wire \malu/_230_ ;
wire \malu/_231_ ;
wire \malu/_232_ ;
wire \malu/_233_ ;
wire \malu/_234_ ;
wire \malu/_235_ ;
wire \malu/_236_ ;
wire \malu/_237_ ;
wire \malu/_238_ ;
wire \malu/_239_ ;
wire \malu/_240_ ;
wire \malu/_241_ ;
wire \malu/_242_ ;
wire \malu/_243_ ;
wire \malu/_244_ ;
wire \malu/_245_ ;
wire \malu/_246_ ;
wire \malu/_247_ ;
wire \malu/_248_ ;
wire \malu/_249_ ;
wire \malu/_250_ ;
wire \malu/_251_ ;
wire \malu/_252_ ;
wire \malu/_253_ ;
wire \malu/_254_ ;
wire \malu/_255_ ;
wire \malu/_256_ ;
wire \malu/_257_ ;
wire \malu/_258_ ;
wire \malu/_259_ ;
wire \malu/_260_ ;
wire \malu/_261_ ;
wire \malu/_262_ ;
wire \malu/_263_ ;
wire \malu/_264_ ;
wire \malu/_265_ ;
wire \malu/_266_ ;
wire \malu/_267_ ;
wire \malu/_268_ ;
wire \malu/_269_ ;
wire \malu/_270_ ;
wire \malu/_271_ ;
wire \malu/_272_ ;
wire \malu/_273_ ;
wire \malu/_274_ ;
wire \malu/_275_ ;
wire \malu/_276_ ;
wire \malu/_277_ ;
wire \malu/_278_ ;
wire \malu/_279_ ;
wire \malu/_280_ ;
wire \malu/_281_ ;
wire \malu/_282_ ;
wire \malu/_283_ ;
wire \malu/_284_ ;
wire \malu/_285_ ;
wire \malu/_286_ ;
wire \malu/_287_ ;
wire \malu/_288_ ;
wire \malu/_289_ ;
wire \malu/_290_ ;
wire \malu/_291_ ;
wire \malu/_292_ ;
wire \malu/_293_ ;
wire \malu/_294_ ;
wire \malu/_295_ ;
wire \malu/_296_ ;
wire \malu/_297_ ;
wire \malu/_298_ ;
wire \malu/_299_ ;
wire \malu/_300_ ;
wire \malu/_301_ ;
wire \malu/_302_ ;
wire \malu/_303_ ;
wire \malu/_304_ ;
wire \malu/_305_ ;
wire \malu/_306_ ;
wire \malu/_307_ ;
wire \malu/adder_result[0] ;
wire \malu/adder_result[10] ;
wire \malu/adder_result[11] ;
wire \malu/adder_result[12] ;
wire \malu/adder_result[13] ;
wire \malu/adder_result[14] ;
wire \malu/adder_result[15] ;
wire \malu/adder_result[16] ;
wire \malu/adder_result[17] ;
wire \malu/adder_result[18] ;
wire \malu/adder_result[19] ;
wire \malu/adder_result[1] ;
wire \malu/adder_result[20] ;
wire \malu/adder_result[21] ;
wire \malu/adder_result[22] ;
wire \malu/adder_result[23] ;
wire \malu/adder_result[24] ;
wire \malu/adder_result[25] ;
wire \malu/adder_result[26] ;
wire \malu/adder_result[27] ;
wire \malu/adder_result[28] ;
wire \malu/adder_result[29] ;
wire \malu/adder_result[2] ;
wire \malu/adder_result[30] ;
wire \malu/adder_result[31] ;
wire \malu/adder_result[3] ;
wire \malu/adder_result[4] ;
wire \malu/adder_result[5] ;
wire \malu/adder_result[6] ;
wire \malu/adder_result[7] ;
wire \malu/adder_result[8] ;
wire \malu/adder_result[9] ;
wire \malu/logic_ctl[0] ;
wire \malu/logic_ctl[1] ;
wire \malu/logic_result[0] ;
wire \malu/logic_result[10] ;
wire \malu/logic_result[11] ;
wire \malu/logic_result[12] ;
wire \malu/logic_result[13] ;
wire \malu/logic_result[14] ;
wire \malu/logic_result[15] ;
wire \malu/logic_result[16] ;
wire \malu/logic_result[17] ;
wire \malu/logic_result[18] ;
wire \malu/logic_result[19] ;
wire \malu/logic_result[1] ;
wire \malu/logic_result[20] ;
wire \malu/logic_result[21] ;
wire \malu/logic_result[22] ;
wire \malu/logic_result[23] ;
wire \malu/logic_result[24] ;
wire \malu/logic_result[25] ;
wire \malu/logic_result[26] ;
wire \malu/logic_result[27] ;
wire \malu/logic_result[28] ;
wire \malu/logic_result[29] ;
wire \malu/logic_result[2] ;
wire \malu/logic_result[30] ;
wire \malu/logic_result[31] ;
wire \malu/logic_result[3] ;
wire \malu/logic_result[4] ;
wire \malu/logic_result[5] ;
wire \malu/logic_result[6] ;
wire \malu/logic_result[7] ;
wire \malu/logic_result[8] ;
wire \malu/logic_result[9] ;
wire \malu/r[0] ;
wire \malu/r[10] ;
wire \malu/r[11] ;
wire \malu/r[12] ;
wire \malu/r[13] ;
wire \malu/r[14] ;
wire \malu/r[15] ;
wire \malu/r[16] ;
wire \malu/r[17] ;
wire \malu/r[18] ;
wire \malu/r[19] ;
wire \malu/r[1] ;
wire \malu/r[20] ;
wire \malu/r[21] ;
wire \malu/r[22] ;
wire \malu/r[23] ;
wire \malu/r[24] ;
wire \malu/r[25] ;
wire \malu/r[26] ;
wire \malu/r[27] ;
wire \malu/r[28] ;
wire \malu/r[29] ;
wire \malu/r[2] ;
wire \malu/r[30] ;
wire \malu/r[31] ;
wire \malu/r[3] ;
wire \malu/r[4] ;
wire \malu/r[5] ;
wire \malu/r[6] ;
wire \malu/r[7] ;
wire \malu/r[8] ;
wire \malu/r[9] ;
wire \malu/shift_ctl[0] ;
wire \malu/shift_ctl[1] ;
wire \malu/shift_result[0] ;
wire \malu/shift_result[10] ;
wire \malu/shift_result[11] ;
wire \malu/shift_result[12] ;
wire \malu/shift_result[13] ;
wire \malu/shift_result[14] ;
wire \malu/shift_result[15] ;
wire \malu/shift_result[16] ;
wire \malu/shift_result[17] ;
wire \malu/shift_result[18] ;
wire \malu/shift_result[19] ;
wire \malu/shift_result[1] ;
wire \malu/shift_result[20] ;
wire \malu/shift_result[21] ;
wire \malu/shift_result[22] ;
wire \malu/shift_result[23] ;
wire \malu/shift_result[24] ;
wire \malu/shift_result[25] ;
wire \malu/shift_result[26] ;
wire \malu/shift_result[27] ;
wire \malu/shift_result[28] ;
wire \malu/shift_result[29] ;
wire \malu/shift_result[2] ;
wire \malu/shift_result[30] ;
wire \malu/shift_result[31] ;
wire \malu/shift_result[3] ;
wire \malu/shift_result[4] ;
wire \malu/shift_result[5] ;
wire \malu/shift_result[6] ;
wire \malu/shift_result[7] ;
wire \malu/shift_result[8] ;
wire \malu/shift_result[9] ;
wire \malu/Adder/_000_ ;
wire \malu/Adder/_001_ ;
wire \malu/Adder/_002_ ;
wire \malu/Adder/_003_ ;
wire \malu/Adder/_004_ ;
wire \malu/Adder/_005_ ;
wire \malu/Adder/_006_ ;
wire \malu/Adder/_007_ ;
wire \malu/Adder/_008_ ;
wire \malu/Adder/_009_ ;
wire \malu/Adder/_010_ ;
wire \malu/Adder/_011_ ;
wire \malu/Adder/_012_ ;
wire \malu/Adder/_013_ ;
wire \malu/Adder/_014_ ;
wire \malu/Adder/_015_ ;
wire \malu/Adder/_016_ ;
wire \malu/Adder/_017_ ;
wire \malu/Adder/_018_ ;
wire \malu/Adder/_019_ ;
wire \malu/Adder/_020_ ;
wire \malu/Adder/_021_ ;
wire \malu/Adder/_022_ ;
wire \malu/Adder/_023_ ;
wire \malu/Adder/_024_ ;
wire \malu/Adder/_025_ ;
wire \malu/Adder/_026_ ;
wire \malu/Adder/_027_ ;
wire \malu/Adder/_028_ ;
wire \malu/Adder/_029_ ;
wire \malu/Adder/_030_ ;
wire \malu/Adder/_031_ ;
wire \malu/Adder/_032_ ;
wire \malu/Adder/_033_ ;
wire \malu/Adder/_034_ ;
wire \malu/Adder/_035_ ;
wire \malu/Adder/_036_ ;
wire \malu/Adder/_037_ ;
wire \malu/Adder/_038_ ;
wire \malu/Adder/_039_ ;
wire \malu/Adder/_040_ ;
wire \malu/Adder/_041_ ;
wire \malu/Adder/_042_ ;
wire \malu/Adder/_043_ ;
wire \malu/Adder/_044_ ;
wire \malu/Adder/_045_ ;
wire \malu/Adder/_046_ ;
wire \malu/Adder/_047_ ;
wire \malu/Adder/_048_ ;
wire \malu/Adder/_049_ ;
wire \malu/Adder/_050_ ;
wire \malu/Adder/_051_ ;
wire \malu/Adder/_052_ ;
wire \malu/Adder/_053_ ;
wire \malu/Adder/_054_ ;
wire \malu/Adder/_055_ ;
wire \malu/Adder/_056_ ;
wire \malu/Adder/_057_ ;
wire \malu/Adder/_058_ ;
wire \malu/Adder/_059_ ;
wire \malu/Adder/_060_ ;
wire \malu/Adder/_061_ ;
wire \malu/Adder/_062_ ;
wire \malu/Adder/_063_ ;
wire \malu/Adder/_064_ ;
wire \malu/Adder/_065_ ;
wire \malu/Adder/_066_ ;
wire \malu/Adder/_067_ ;
wire \malu/Adder/_068_ ;
wire \malu/Adder/_069_ ;
wire \malu/Adder/_070_ ;
wire \malu/Adder/_071_ ;
wire \malu/Adder/_072_ ;
wire \malu/Adder/_073_ ;
wire \malu/Adder/_074_ ;
wire \malu/Adder/_075_ ;
wire \malu/Adder/_076_ ;
wire \malu/Adder/_077_ ;
wire \malu/Adder/_078_ ;
wire \malu/Adder/_079_ ;
wire \malu/Adder/_080_ ;
wire \malu/Adder/_081_ ;
wire \malu/Adder/_082_ ;
wire \malu/Adder/_083_ ;
wire \malu/Adder/_084_ ;
wire \malu/Adder/_085_ ;
wire \malu/Adder/_086_ ;
wire \malu/Adder/_087_ ;
wire \malu/Adder/_088_ ;
wire \malu/Adder/_089_ ;
wire \malu/Adder/_090_ ;
wire \malu/Adder/_091_ ;
wire \malu/Adder/_092_ ;
wire \malu/Adder/_093_ ;
wire \malu/Adder/_094_ ;
wire \malu/Adder/_095_ ;
wire \malu/Adder/_096_ ;
wire \malu/Adder/_097_ ;
wire \malu/Adder/_098_ ;
wire \malu/Adder/_099_ ;
wire \malu/Adder/_100_ ;
wire \malu/Adder/_101_ ;
wire \malu/Adder/_102_ ;
wire \malu/Adder/_103_ ;
wire \malu/Adder/_104_ ;
wire \malu/Adder/_105_ ;
wire \malu/Adder/_106_ ;
wire \malu/Adder/_107_ ;
wire \malu/Adder/_108_ ;
wire \malu/Adder/_109_ ;
wire \malu/Adder/_110_ ;
wire \malu/Adder/_111_ ;
wire \malu/Adder/_112_ ;
wire \malu/Adder/_113_ ;
wire \malu/Adder/_114_ ;
wire \malu/Adder/_115_ ;
wire \malu/Adder/_116_ ;
wire \malu/Adder/_117_ ;
wire \malu/Adder/_118_ ;
wire \malu/Adder/_119_ ;
wire \malu/Adder/_120_ ;
wire \malu/Adder/_121_ ;
wire \malu/Adder/_122_ ;
wire \malu/Adder/_123_ ;
wire \malu/Adder/_124_ ;
wire \malu/Adder/_125_ ;
wire \malu/Adder/_126_ ;
wire \malu/Adder/_127_ ;
wire \malu/Adder/_128_ ;
wire \malu/Adder/_129_ ;
wire \malu/Adder/_130_ ;
wire \malu/Adder/_131_ ;
wire \malu/Adder/_132_ ;
wire \malu/Adder/_133_ ;
wire \malu/Adder/_134_ ;
wire \malu/Adder/_135_ ;
wire \malu/Adder/_136_ ;
wire \malu/Adder/_137_ ;
wire \malu/Adder/_138_ ;
wire \malu/Adder/_139_ ;
wire \malu/Adder/_140_ ;
wire \malu/Adder/_141_ ;
wire \malu/Adder/_142_ ;
wire \malu/Adder/_143_ ;
wire \malu/Adder/_144_ ;
wire \malu/Adder/_145_ ;
wire \malu/Adder/_146_ ;
wire \malu/Adder/_147_ ;
wire \malu/Adder/_148_ ;
wire \malu/Adder/_149_ ;
wire \malu/Adder/_150_ ;
wire \malu/Adder/_151_ ;
wire \malu/Adder/_152_ ;
wire \malu/Adder/_153_ ;
wire \malu/Adder/_154_ ;
wire \malu/Adder/_155_ ;
wire \malu/Adder/_156_ ;
wire \malu/Adder/_157_ ;
wire \malu/Adder/_158_ ;
wire \malu/Adder/_159_ ;
wire \malu/Adder/_160_ ;
wire \malu/Adder/_161_ ;
wire \malu/Adder/_162_ ;
wire \malu/Adder/_163_ ;
wire \malu/Adder/_164_ ;
wire \malu/Adder/_165_ ;
wire \malu/Adder/_166_ ;
wire \malu/Adder/_167_ ;
wire \malu/Adder/_168_ ;
wire \malu/Adder/_169_ ;
wire \malu/Adder/_170_ ;
wire \malu/Adder/_171_ ;
wire \malu/Adder/_172_ ;
wire \malu/Adder/_173_ ;
wire \malu/Adder/_174_ ;
wire \malu/Adder/_175_ ;
wire \malu/Adder/_176_ ;
wire \malu/Adder/_177_ ;
wire \malu/Adder/_178_ ;
wire \malu/Adder/_179_ ;
wire \malu/Adder/_180_ ;
wire \malu/Adder/_181_ ;
wire \malu/Adder/_182_ ;
wire \malu/Adder/_183_ ;
wire \malu/Adder/_184_ ;
wire \malu/Adder/_185_ ;
wire \malu/Adder/_186_ ;
wire \malu/Adder/_187_ ;
wire \malu/Adder/_188_ ;
wire \malu/Adder/_189_ ;
wire \malu/Adder/_190_ ;
wire \malu/Adder/_191_ ;
wire \malu/Adder/_192_ ;
wire \malu/Adder/_193_ ;
wire \malu/Adder/_194_ ;
wire \malu/Adder/_195_ ;
wire \malu/Adder/_196_ ;
wire \malu/Adder/_197_ ;
wire \malu/Adder/_198_ ;
wire \malu/Adder/_199_ ;
wire \malu/Adder/_200_ ;
wire \malu/Adder/_201_ ;
wire \malu/Adder/_202_ ;
wire \malu/Adder/_203_ ;
wire \malu/Adder/_204_ ;
wire \malu/Adder/_205_ ;
wire \malu/Adder/_206_ ;
wire \malu/Adder/_207_ ;
wire \malu/Adder/_208_ ;
wire \malu/Adder/_209_ ;
wire \malu/Adder/_210_ ;
wire \malu/Adder/_211_ ;
wire \malu/Adder/_212_ ;
wire \malu/Adder/_213_ ;
wire \malu/Adder/_214_ ;
wire \malu/Adder/_215_ ;
wire \malu/Adder/_216_ ;
wire \malu/Adder/_217_ ;
wire \malu/Adder/_218_ ;
wire \malu/Adder/_219_ ;
wire \malu/Adder/_220_ ;
wire \malu/Adder/_221_ ;
wire \malu/Adder/_222_ ;
wire \malu/Adder/_223_ ;
wire \malu/Adder/_224_ ;
wire \malu/Adder/_225_ ;
wire \malu/Adder/_226_ ;
wire \malu/Adder/_227_ ;
wire \malu/Adder/_228_ ;
wire \malu/Adder/_229_ ;
wire \malu/Adder/_230_ ;
wire \malu/Adder/_231_ ;
wire \malu/Adder/_232_ ;
wire \malu/Adder/_233_ ;
wire \malu/Adder/_234_ ;
wire \malu/Adder/_235_ ;
wire \malu/Adder/_236_ ;
wire \malu/Adder/_237_ ;
wire \malu/Adder/_238_ ;
wire \malu/Adder/_239_ ;
wire \malu/Adder/_240_ ;
wire \malu/Adder/_241_ ;
wire \malu/Adder/_242_ ;
wire \malu/Adder/_243_ ;
wire \malu/Adder/_244_ ;
wire \malu/Adder/_245_ ;
wire \malu/Adder/_246_ ;
wire \malu/Adder/_247_ ;
wire \malu/Adder/_248_ ;
wire \malu/Adder/_249_ ;
wire \malu/Adder/_250_ ;
wire \malu/Adder/_251_ ;
wire \malu/Adder/_252_ ;
wire \malu/Adder/_253_ ;
wire \malu/Adder/_254_ ;
wire \malu/Adder/_255_ ;
wire \malu/Adder/_256_ ;
wire \malu/Adder/_257_ ;
wire \malu/Adder/_258_ ;
wire \malu/Adder/_259_ ;
wire \malu/Adder/_260_ ;
wire \malu/Adder/_261_ ;
wire \malu/Adder/_262_ ;
wire \malu/Adder/_263_ ;
wire \malu/Adder/_264_ ;
wire \malu/Adder/_265_ ;
wire \malu/Adder/_266_ ;
wire \malu/Adder/_267_ ;
wire \malu/Adder/_268_ ;
wire \malu/Adder/_269_ ;
wire \malu/Adder/_270_ ;
wire \malu/Adder/_271_ ;
wire \malu/Adder/_272_ ;
wire \malu/Adder/_273_ ;
wire \malu/Adder/_274_ ;
wire \malu/Adder/_275_ ;
wire \malu/Adder/_276_ ;
wire \malu/Adder/_277_ ;
wire \malu/Adder/_278_ ;
wire \malu/Adder/_279_ ;
wire \malu/Adder/_280_ ;
wire \malu/Adder/_281_ ;
wire \malu/Adder/_282_ ;
wire \malu/Adder/_283_ ;
wire \malu/Adder/_284_ ;
wire \malu/Adder/_285_ ;
wire \malu/Adder/_286_ ;
wire \malu/Adder/_287_ ;
wire \malu/Adder/_288_ ;
wire \malu/Adder/_289_ ;
wire \malu/Adder/_290_ ;
wire \malu/Adder/_291_ ;
wire \malu/Adder/_292_ ;
wire \malu/Adder/_293_ ;
wire \malu/Adder/_294_ ;
wire \malu/Adder/_295_ ;
wire \malu/Adder/_296_ ;
wire \malu/Adder/_297_ ;
wire \malu/Adder/_298_ ;
wire \malu/Adder/_299_ ;
wire \malu/Adder/_300_ ;
wire \malu/Adder/_301_ ;
wire \malu/Adder/_302_ ;
wire \malu/Adder/_303_ ;
wire \malu/Adder/_304_ ;
wire \malu/Adder/_305_ ;
wire \malu/Adder/_306_ ;
wire \malu/Adder/_307_ ;
wire \malu/Adder/_308_ ;
wire \malu/Adder/_309_ ;
wire \malu/Adder/_310_ ;
wire \malu/Adder/_311_ ;
wire \malu/Adder/_312_ ;
wire \malu/Adder/_313_ ;
wire \malu/Adder/_314_ ;
wire \malu/Adder/_315_ ;
wire \malu/Adder/_316_ ;
wire \malu/Adder/_317_ ;
wire \malu/Adder/_318_ ;
wire \malu/Adder/_319_ ;
wire \malu/Adder/_320_ ;
wire \malu/Adder/_321_ ;
wire \malu/Adder/_322_ ;
wire \malu/Adder/_323_ ;
wire \malu/Logic/_000_ ;
wire \malu/Logic/_001_ ;
wire \malu/Logic/_002_ ;
wire \malu/Logic/_003_ ;
wire \malu/Logic/_004_ ;
wire \malu/Logic/_005_ ;
wire \malu/Logic/_006_ ;
wire \malu/Logic/_007_ ;
wire \malu/Logic/_008_ ;
wire \malu/Logic/_009_ ;
wire \malu/Logic/_010_ ;
wire \malu/Logic/_011_ ;
wire \malu/Logic/_012_ ;
wire \malu/Logic/_013_ ;
wire \malu/Logic/_014_ ;
wire \malu/Logic/_015_ ;
wire \malu/Logic/_016_ ;
wire \malu/Logic/_017_ ;
wire \malu/Logic/_018_ ;
wire \malu/Logic/_019_ ;
wire \malu/Logic/_020_ ;
wire \malu/Logic/_021_ ;
wire \malu/Logic/_022_ ;
wire \malu/Logic/_023_ ;
wire \malu/Logic/_024_ ;
wire \malu/Logic/_025_ ;
wire \malu/Logic/_026_ ;
wire \malu/Logic/_027_ ;
wire \malu/Logic/_028_ ;
wire \malu/Logic/_029_ ;
wire \malu/Logic/_030_ ;
wire \malu/Logic/_031_ ;
wire \malu/Logic/_032_ ;
wire \malu/Logic/_033_ ;
wire \malu/Logic/_034_ ;
wire \malu/Logic/_035_ ;
wire \malu/Logic/_036_ ;
wire \malu/Logic/_037_ ;
wire \malu/Logic/_038_ ;
wire \malu/Logic/_039_ ;
wire \malu/Logic/_040_ ;
wire \malu/Logic/_041_ ;
wire \malu/Logic/_042_ ;
wire \malu/Logic/_043_ ;
wire \malu/Logic/_044_ ;
wire \malu/Logic/_045_ ;
wire \malu/Logic/_046_ ;
wire \malu/Logic/_047_ ;
wire \malu/Logic/_048_ ;
wire \malu/Logic/_049_ ;
wire \malu/Logic/_050_ ;
wire \malu/Logic/_051_ ;
wire \malu/Logic/_052_ ;
wire \malu/Logic/_053_ ;
wire \malu/Logic/_054_ ;
wire \malu/Logic/_055_ ;
wire \malu/Logic/_056_ ;
wire \malu/Logic/_057_ ;
wire \malu/Logic/_058_ ;
wire \malu/Logic/_059_ ;
wire \malu/Logic/_060_ ;
wire \malu/Logic/_061_ ;
wire \malu/Logic/_062_ ;
wire \malu/Logic/_063_ ;
wire \malu/Logic/_064_ ;
wire \malu/Logic/_065_ ;
wire \malu/Logic/_066_ ;
wire \malu/Logic/_067_ ;
wire \malu/Logic/_068_ ;
wire \malu/Logic/_069_ ;
wire \malu/Logic/_070_ ;
wire \malu/Logic/_071_ ;
wire \malu/Logic/_072_ ;
wire \malu/Logic/_073_ ;
wire \malu/Logic/_074_ ;
wire \malu/Logic/_075_ ;
wire \malu/Logic/_076_ ;
wire \malu/Logic/_077_ ;
wire \malu/Logic/_078_ ;
wire \malu/Logic/_079_ ;
wire \malu/Logic/_080_ ;
wire \malu/Logic/_081_ ;
wire \malu/Logic/_082_ ;
wire \malu/Logic/_083_ ;
wire \malu/Logic/_084_ ;
wire \malu/Logic/_085_ ;
wire \malu/Logic/_086_ ;
wire \malu/Logic/_087_ ;
wire \malu/Logic/_088_ ;
wire \malu/Logic/_089_ ;
wire \malu/Logic/_090_ ;
wire \malu/Logic/_091_ ;
wire \malu/Logic/_092_ ;
wire \malu/Logic/_093_ ;
wire \malu/Logic/_094_ ;
wire \malu/Logic/_095_ ;
wire \malu/Logic/_096_ ;
wire \malu/Logic/_097_ ;
wire \malu/Logic/_098_ ;
wire \malu/Logic/_099_ ;
wire \malu/Logic/_100_ ;
wire \malu/Logic/_101_ ;
wire \malu/Logic/_102_ ;
wire \malu/Logic/_103_ ;
wire \malu/Logic/_104_ ;
wire \malu/Logic/_105_ ;
wire \malu/Logic/_106_ ;
wire \malu/Logic/_107_ ;
wire \malu/Logic/_108_ ;
wire \malu/Logic/_109_ ;
wire \malu/Logic/_110_ ;
wire \malu/Logic/_111_ ;
wire \malu/Logic/_112_ ;
wire \malu/Logic/_113_ ;
wire \malu/Logic/_114_ ;
wire \malu/Logic/_115_ ;
wire \malu/Logic/_116_ ;
wire \malu/Logic/_117_ ;
wire \malu/Logic/_118_ ;
wire \malu/Logic/_119_ ;
wire \malu/Logic/_120_ ;
wire \malu/Logic/_121_ ;
wire \malu/Logic/_122_ ;
wire \malu/Logic/_123_ ;
wire \malu/Logic/_124_ ;
wire \malu/Logic/_125_ ;
wire \malu/Logic/_126_ ;
wire \malu/Logic/_127_ ;
wire \malu/Logic/_128_ ;
wire \malu/Logic/_129_ ;
wire \malu/Logic/_130_ ;
wire \malu/Logic/_131_ ;
wire \malu/Logic/_132_ ;
wire \malu/Logic/_133_ ;
wire \malu/Logic/_134_ ;
wire \malu/Logic/_135_ ;
wire \malu/Logic/_136_ ;
wire \malu/Logic/_137_ ;
wire \malu/Logic/_138_ ;
wire \malu/Logic/_139_ ;
wire \malu/Logic/_140_ ;
wire \malu/Logic/_141_ ;
wire \malu/Logic/_142_ ;
wire \malu/Logic/_143_ ;
wire \malu/Logic/_144_ ;
wire \malu/Logic/_145_ ;
wire \malu/Logic/_146_ ;
wire \malu/Logic/_147_ ;
wire \malu/Logic/_148_ ;
wire \malu/Logic/_149_ ;
wire \malu/Logic/_150_ ;
wire \malu/Logic/_151_ ;
wire \malu/Logic/_152_ ;
wire \malu/Logic/_153_ ;
wire \malu/Logic/_154_ ;
wire \malu/Logic/_155_ ;
wire \malu/Logic/_156_ ;
wire \malu/Logic/_157_ ;
wire \malu/Logic/_158_ ;
wire \malu/Logic/_159_ ;
wire \malu/Logic/_160_ ;
wire \malu/Logic/_161_ ;
wire \malu/Logic/_162_ ;
wire \malu/Logic/_163_ ;
wire \malu/Logic/_164_ ;
wire \malu/Logic/_165_ ;
wire \malu/Logic/_166_ ;
wire \malu/Logic/_167_ ;
wire \malu/Logic/_168_ ;
wire \malu/Logic/_169_ ;
wire \malu/Logic/_170_ ;
wire \malu/Logic/_171_ ;
wire \malu/Logic/_172_ ;
wire \malu/Logic/_173_ ;
wire \malu/Logic/_174_ ;
wire \malu/Logic/_175_ ;
wire \malu/Logic/_176_ ;
wire \malu/Logic/_177_ ;
wire \malu/Logic/_178_ ;
wire \malu/Logic/_179_ ;
wire \malu/Logic/_180_ ;
wire \malu/Logic/_181_ ;
wire \malu/Logic/_182_ ;
wire \malu/Logic/_183_ ;
wire \malu/Logic/_184_ ;
wire \malu/Logic/_185_ ;
wire \malu/Logic/_186_ ;
wire \malu/Logic/_187_ ;
wire \malu/Logic/_188_ ;
wire \malu/Logic/_189_ ;
wire \malu/Logic/_190_ ;
wire \malu/Logic/_191_ ;
wire \malu/Logic/_192_ ;
wire \malu/Logic/_193_ ;
wire \malu/Logic/_194_ ;
wire \malu/Logic/_195_ ;
wire \malu/Logic/_196_ ;
wire \malu/Logic/_197_ ;
wire \malu/Logic/_198_ ;
wire \malu/Logic/_199_ ;
wire \malu/Logic/_200_ ;
wire \malu/Logic/_201_ ;
wire \malu/Shift/_0000_ ;
wire \malu/Shift/_0001_ ;
wire \malu/Shift/_0002_ ;
wire \malu/Shift/_0003_ ;
wire \malu/Shift/_0004_ ;
wire \malu/Shift/_0005_ ;
wire \malu/Shift/_0006_ ;
wire \malu/Shift/_0007_ ;
wire \malu/Shift/_0008_ ;
wire \malu/Shift/_0009_ ;
wire \malu/Shift/_0010_ ;
wire \malu/Shift/_0011_ ;
wire \malu/Shift/_0012_ ;
wire \malu/Shift/_0013_ ;
wire \malu/Shift/_0014_ ;
wire \malu/Shift/_0015_ ;
wire \malu/Shift/_0016_ ;
wire \malu/Shift/_0017_ ;
wire \malu/Shift/_0018_ ;
wire \malu/Shift/_0019_ ;
wire \malu/Shift/_0020_ ;
wire \malu/Shift/_0021_ ;
wire \malu/Shift/_0022_ ;
wire \malu/Shift/_0023_ ;
wire \malu/Shift/_0024_ ;
wire \malu/Shift/_0025_ ;
wire \malu/Shift/_0026_ ;
wire \malu/Shift/_0027_ ;
wire \malu/Shift/_0028_ ;
wire \malu/Shift/_0029_ ;
wire \malu/Shift/_0030_ ;
wire \malu/Shift/_0031_ ;
wire \malu/Shift/_0032_ ;
wire \malu/Shift/_0033_ ;
wire \malu/Shift/_0034_ ;
wire \malu/Shift/_0035_ ;
wire \malu/Shift/_0036_ ;
wire \malu/Shift/_0037_ ;
wire \malu/Shift/_0038_ ;
wire \malu/Shift/_0039_ ;
wire \malu/Shift/_0040_ ;
wire \malu/Shift/_0041_ ;
wire \malu/Shift/_0042_ ;
wire \malu/Shift/_0043_ ;
wire \malu/Shift/_0044_ ;
wire \malu/Shift/_0045_ ;
wire \malu/Shift/_0046_ ;
wire \malu/Shift/_0047_ ;
wire \malu/Shift/_0048_ ;
wire \malu/Shift/_0049_ ;
wire \malu/Shift/_0050_ ;
wire \malu/Shift/_0051_ ;
wire \malu/Shift/_0052_ ;
wire \malu/Shift/_0053_ ;
wire \malu/Shift/_0054_ ;
wire \malu/Shift/_0055_ ;
wire \malu/Shift/_0056_ ;
wire \malu/Shift/_0057_ ;
wire \malu/Shift/_0058_ ;
wire \malu/Shift/_0059_ ;
wire \malu/Shift/_0060_ ;
wire \malu/Shift/_0061_ ;
wire \malu/Shift/_0062_ ;
wire \malu/Shift/_0063_ ;
wire \malu/Shift/_0064_ ;
wire \malu/Shift/_0065_ ;
wire \malu/Shift/_0066_ ;
wire \malu/Shift/_0067_ ;
wire \malu/Shift/_0068_ ;
wire \malu/Shift/_0069_ ;
wire \malu/Shift/_0070_ ;
wire \malu/Shift/_0071_ ;
wire \malu/Shift/_0072_ ;
wire \malu/Shift/_0073_ ;
wire \malu/Shift/_0074_ ;
wire \malu/Shift/_0075_ ;
wire \malu/Shift/_0076_ ;
wire \malu/Shift/_0077_ ;
wire \malu/Shift/_0078_ ;
wire \malu/Shift/_0079_ ;
wire \malu/Shift/_0080_ ;
wire \malu/Shift/_0081_ ;
wire \malu/Shift/_0082_ ;
wire \malu/Shift/_0083_ ;
wire \malu/Shift/_0084_ ;
wire \malu/Shift/_0085_ ;
wire \malu/Shift/_0086_ ;
wire \malu/Shift/_0087_ ;
wire \malu/Shift/_0088_ ;
wire \malu/Shift/_0089_ ;
wire \malu/Shift/_0090_ ;
wire \malu/Shift/_0091_ ;
wire \malu/Shift/_0092_ ;
wire \malu/Shift/_0093_ ;
wire \malu/Shift/_0094_ ;
wire \malu/Shift/_0095_ ;
wire \malu/Shift/_0096_ ;
wire \malu/Shift/_0097_ ;
wire \malu/Shift/_0098_ ;
wire \malu/Shift/_0099_ ;
wire \malu/Shift/_0100_ ;
wire \malu/Shift/_0101_ ;
wire \malu/Shift/_0102_ ;
wire \malu/Shift/_0103_ ;
wire \malu/Shift/_0104_ ;
wire \malu/Shift/_0105_ ;
wire \malu/Shift/_0106_ ;
wire \malu/Shift/_0107_ ;
wire \malu/Shift/_0108_ ;
wire \malu/Shift/_0109_ ;
wire \malu/Shift/_0110_ ;
wire \malu/Shift/_0111_ ;
wire \malu/Shift/_0112_ ;
wire \malu/Shift/_0113_ ;
wire \malu/Shift/_0114_ ;
wire \malu/Shift/_0115_ ;
wire \malu/Shift/_0116_ ;
wire \malu/Shift/_0117_ ;
wire \malu/Shift/_0118_ ;
wire \malu/Shift/_0119_ ;
wire \malu/Shift/_0120_ ;
wire \malu/Shift/_0121_ ;
wire \malu/Shift/_0122_ ;
wire \malu/Shift/_0123_ ;
wire \malu/Shift/_0124_ ;
wire \malu/Shift/_0125_ ;
wire \malu/Shift/_0126_ ;
wire \malu/Shift/_0127_ ;
wire \malu/Shift/_0128_ ;
wire \malu/Shift/_0129_ ;
wire \malu/Shift/_0130_ ;
wire \malu/Shift/_0131_ ;
wire \malu/Shift/_0132_ ;
wire \malu/Shift/_0133_ ;
wire \malu/Shift/_0134_ ;
wire \malu/Shift/_0135_ ;
wire \malu/Shift/_0136_ ;
wire \malu/Shift/_0137_ ;
wire \malu/Shift/_0138_ ;
wire \malu/Shift/_0139_ ;
wire \malu/Shift/_0140_ ;
wire \malu/Shift/_0141_ ;
wire \malu/Shift/_0142_ ;
wire \malu/Shift/_0143_ ;
wire \malu/Shift/_0144_ ;
wire \malu/Shift/_0145_ ;
wire \malu/Shift/_0146_ ;
wire \malu/Shift/_0147_ ;
wire \malu/Shift/_0148_ ;
wire \malu/Shift/_0149_ ;
wire \malu/Shift/_0150_ ;
wire \malu/Shift/_0151_ ;
wire \malu/Shift/_0152_ ;
wire \malu/Shift/_0153_ ;
wire \malu/Shift/_0154_ ;
wire \malu/Shift/_0155_ ;
wire \malu/Shift/_0156_ ;
wire \malu/Shift/_0157_ ;
wire \malu/Shift/_0158_ ;
wire \malu/Shift/_0159_ ;
wire \malu/Shift/_0160_ ;
wire \malu/Shift/_0161_ ;
wire \malu/Shift/_0162_ ;
wire \malu/Shift/_0163_ ;
wire \malu/Shift/_0164_ ;
wire \malu/Shift/_0165_ ;
wire \malu/Shift/_0166_ ;
wire \malu/Shift/_0167_ ;
wire \malu/Shift/_0168_ ;
wire \malu/Shift/_0169_ ;
wire \malu/Shift/_0170_ ;
wire \malu/Shift/_0171_ ;
wire \malu/Shift/_0172_ ;
wire \malu/Shift/_0173_ ;
wire \malu/Shift/_0174_ ;
wire \malu/Shift/_0175_ ;
wire \malu/Shift/_0176_ ;
wire \malu/Shift/_0177_ ;
wire \malu/Shift/_0178_ ;
wire \malu/Shift/_0179_ ;
wire \malu/Shift/_0180_ ;
wire \malu/Shift/_0181_ ;
wire \malu/Shift/_0182_ ;
wire \malu/Shift/_0183_ ;
wire \malu/Shift/_0184_ ;
wire \malu/Shift/_0185_ ;
wire \malu/Shift/_0186_ ;
wire \malu/Shift/_0187_ ;
wire \malu/Shift/_0188_ ;
wire \malu/Shift/_0189_ ;
wire \malu/Shift/_0190_ ;
wire \malu/Shift/_0191_ ;
wire \malu/Shift/_0192_ ;
wire \malu/Shift/_0193_ ;
wire \malu/Shift/_0194_ ;
wire \malu/Shift/_0195_ ;
wire \malu/Shift/_0196_ ;
wire \malu/Shift/_0197_ ;
wire \malu/Shift/_0198_ ;
wire \malu/Shift/_0199_ ;
wire \malu/Shift/_0200_ ;
wire \malu/Shift/_0201_ ;
wire \malu/Shift/_0202_ ;
wire \malu/Shift/_0203_ ;
wire \malu/Shift/_0204_ ;
wire \malu/Shift/_0205_ ;
wire \malu/Shift/_0206_ ;
wire \malu/Shift/_0207_ ;
wire \malu/Shift/_0208_ ;
wire \malu/Shift/_0209_ ;
wire \malu/Shift/_0210_ ;
wire \malu/Shift/_0211_ ;
wire \malu/Shift/_0212_ ;
wire \malu/Shift/_0213_ ;
wire \malu/Shift/_0214_ ;
wire \malu/Shift/_0215_ ;
wire \malu/Shift/_0216_ ;
wire \malu/Shift/_0217_ ;
wire \malu/Shift/_0218_ ;
wire \malu/Shift/_0219_ ;
wire \malu/Shift/_0220_ ;
wire \malu/Shift/_0221_ ;
wire \malu/Shift/_0222_ ;
wire \malu/Shift/_0223_ ;
wire \malu/Shift/_0224_ ;
wire \malu/Shift/_0225_ ;
wire \malu/Shift/_0226_ ;
wire \malu/Shift/_0227_ ;
wire \malu/Shift/_0228_ ;
wire \malu/Shift/_0229_ ;
wire \malu/Shift/_0230_ ;
wire \malu/Shift/_0231_ ;
wire \malu/Shift/_0232_ ;
wire \malu/Shift/_0233_ ;
wire \malu/Shift/_0234_ ;
wire \malu/Shift/_0235_ ;
wire \malu/Shift/_0236_ ;
wire \malu/Shift/_0237_ ;
wire \malu/Shift/_0238_ ;
wire \malu/Shift/_0239_ ;
wire \malu/Shift/_0240_ ;
wire \malu/Shift/_0241_ ;
wire \malu/Shift/_0242_ ;
wire \malu/Shift/_0243_ ;
wire \malu/Shift/_0244_ ;
wire \malu/Shift/_0245_ ;
wire \malu/Shift/_0246_ ;
wire \malu/Shift/_0247_ ;
wire \malu/Shift/_0248_ ;
wire \malu/Shift/_0249_ ;
wire \malu/Shift/_0250_ ;
wire \malu/Shift/_0251_ ;
wire \malu/Shift/_0252_ ;
wire \malu/Shift/_0253_ ;
wire \malu/Shift/_0254_ ;
wire \malu/Shift/_0255_ ;
wire \malu/Shift/_0256_ ;
wire \malu/Shift/_0257_ ;
wire \malu/Shift/_0258_ ;
wire \malu/Shift/_0259_ ;
wire \malu/Shift/_0260_ ;
wire \malu/Shift/_0261_ ;
wire \malu/Shift/_0262_ ;
wire \malu/Shift/_0263_ ;
wire \malu/Shift/_0264_ ;
wire \malu/Shift/_0265_ ;
wire \malu/Shift/_0266_ ;
wire \malu/Shift/_0267_ ;
wire \malu/Shift/_0268_ ;
wire \malu/Shift/_0269_ ;
wire \malu/Shift/_0270_ ;
wire \malu/Shift/_0271_ ;
wire \malu/Shift/_0272_ ;
wire \malu/Shift/_0273_ ;
wire \malu/Shift/_0274_ ;
wire \malu/Shift/_0275_ ;
wire \malu/Shift/_0276_ ;
wire \malu/Shift/_0277_ ;
wire \malu/Shift/_0278_ ;
wire \malu/Shift/_0279_ ;
wire \malu/Shift/_0280_ ;
wire \malu/Shift/_0281_ ;
wire \malu/Shift/_0282_ ;
wire \malu/Shift/_0283_ ;
wire \malu/Shift/_0284_ ;
wire \malu/Shift/_0285_ ;
wire \malu/Shift/_0286_ ;
wire \malu/Shift/_0287_ ;
wire \malu/Shift/_0288_ ;
wire \malu/Shift/_0289_ ;
wire \malu/Shift/_0290_ ;
wire \malu/Shift/_0291_ ;
wire \malu/Shift/_0292_ ;
wire \malu/Shift/_0293_ ;
wire \malu/Shift/_0294_ ;
wire \malu/Shift/_0295_ ;
wire \malu/Shift/_0296_ ;
wire \malu/Shift/_0297_ ;
wire \malu/Shift/_0298_ ;
wire \malu/Shift/_0299_ ;
wire \malu/Shift/_0300_ ;
wire \malu/Shift/_0301_ ;
wire \malu/Shift/_0302_ ;
wire \malu/Shift/_0303_ ;
wire \malu/Shift/_0304_ ;
wire \malu/Shift/_0305_ ;
wire \malu/Shift/_0306_ ;
wire \malu/Shift/_0307_ ;
wire \malu/Shift/_0308_ ;
wire \malu/Shift/_0309_ ;
wire \malu/Shift/_0310_ ;
wire \malu/Shift/_0311_ ;
wire \malu/Shift/_0312_ ;
wire \malu/Shift/_0313_ ;
wire \malu/Shift/_0314_ ;
wire \malu/Shift/_0315_ ;
wire \malu/Shift/_0316_ ;
wire \malu/Shift/_0317_ ;
wire \malu/Shift/_0318_ ;
wire \malu/Shift/_0319_ ;
wire \malu/Shift/_0320_ ;
wire \malu/Shift/_0321_ ;
wire \malu/Shift/_0322_ ;
wire \malu/Shift/_0323_ ;
wire \malu/Shift/_0324_ ;
wire \malu/Shift/_0325_ ;
wire \malu/Shift/_0326_ ;
wire \malu/Shift/_0327_ ;
wire \malu/Shift/_0328_ ;
wire \malu/Shift/_0329_ ;
wire \malu/Shift/_0330_ ;
wire \malu/Shift/_0331_ ;
wire \malu/Shift/_0332_ ;
wire \malu/Shift/_0333_ ;
wire \malu/Shift/_0334_ ;
wire \malu/Shift/_0335_ ;
wire \malu/Shift/_0336_ ;
wire \malu/Shift/_0337_ ;
wire \malu/Shift/_0338_ ;
wire \malu/Shift/_0339_ ;
wire \malu/Shift/_0340_ ;
wire \malu/Shift/_0341_ ;
wire \malu/Shift/_0342_ ;
wire \malu/Shift/_0343_ ;
wire \malu/Shift/_0344_ ;
wire \malu/Shift/_0345_ ;
wire \malu/Shift/_0346_ ;
wire \malu/Shift/_0347_ ;
wire \malu/Shift/_0348_ ;
wire \malu/Shift/_0349_ ;
wire \malu/Shift/_0350_ ;
wire \malu/Shift/_0351_ ;
wire \malu/Shift/_0352_ ;
wire \malu/Shift/_0353_ ;
wire \malu/Shift/_0354_ ;
wire \malu/Shift/_0355_ ;
wire \malu/Shift/_0356_ ;
wire \malu/Shift/_0357_ ;
wire \malu/Shift/_0358_ ;
wire \malu/Shift/_0359_ ;
wire \malu/Shift/_0360_ ;
wire \malu/Shift/_0361_ ;
wire \malu/Shift/_0362_ ;
wire \malu/Shift/_0363_ ;
wire \malu/Shift/_0364_ ;
wire \malu/Shift/_0365_ ;
wire \malu/Shift/_0366_ ;
wire \malu/Shift/_0367_ ;
wire \malu/Shift/_0368_ ;
wire \malu/Shift/_0369_ ;
wire \malu/Shift/_0370_ ;
wire \malu/Shift/_0371_ ;
wire \malu/Shift/_0372_ ;
wire \malu/Shift/_0373_ ;
wire \malu/Shift/_0374_ ;
wire \malu/Shift/_0375_ ;
wire \malu/Shift/_0376_ ;
wire \malu/Shift/_0377_ ;
wire \malu/Shift/_0378_ ;
wire \malu/Shift/_0379_ ;
wire \malu/Shift/_0380_ ;
wire \malu/Shift/_0381_ ;
wire \malu/Shift/_0382_ ;
wire \malu/Shift/_0383_ ;
wire \malu/Shift/_0384_ ;
wire \malu/Shift/_0385_ ;
wire \malu/Shift/_0386_ ;
wire \malu/Shift/_0387_ ;
wire \malu/Shift/_0388_ ;
wire \malu/Shift/_0389_ ;
wire \malu/Shift/_0390_ ;
wire \malu/Shift/_0391_ ;
wire \malu/Shift/_0392_ ;
wire \malu/Shift/_0393_ ;
wire \malu/Shift/_0394_ ;
wire \malu/Shift/_0395_ ;
wire \malu/Shift/_0396_ ;
wire \malu/Shift/_0397_ ;
wire \malu/Shift/_0398_ ;
wire \malu/Shift/_0399_ ;
wire \malu/Shift/_0400_ ;
wire \malu/Shift/_0401_ ;
wire \malu/Shift/_0402_ ;
wire \malu/Shift/_0403_ ;
wire \malu/Shift/_0404_ ;
wire \malu/Shift/_0405_ ;
wire \malu/Shift/_0406_ ;
wire \malu/Shift/_0407_ ;
wire \malu/Shift/_0408_ ;
wire \malu/Shift/_0409_ ;
wire \malu/Shift/_0410_ ;
wire \malu/Shift/_0411_ ;
wire \malu/Shift/_0412_ ;
wire \malu/Shift/_0413_ ;
wire \malu/Shift/_0414_ ;
wire \malu/Shift/_0415_ ;
wire \malu/Shift/_0416_ ;
wire \malu/Shift/_0417_ ;
wire \malu/Shift/_0418_ ;
wire \malu/Shift/_0419_ ;
wire \malu/Shift/_0420_ ;
wire \malu/Shift/_0421_ ;
wire \malu/Shift/_0422_ ;
wire \malu/Shift/_0423_ ;
wire \malu/Shift/_0424_ ;
wire \malu/Shift/_0425_ ;
wire \malu/Shift/_0426_ ;
wire \malu/Shift/_0427_ ;
wire \malu/Shift/_0428_ ;
wire \malu/Shift/_0429_ ;
wire \malu/Shift/_0430_ ;
wire \malu/Shift/_0431_ ;
wire \malu/Shift/_0432_ ;
wire \malu/Shift/_0433_ ;
wire \malu/Shift/_0434_ ;
wire \malu/Shift/_0435_ ;
wire \malu/Shift/_0436_ ;
wire \malu/Shift/_0437_ ;
wire \malu/Shift/_0438_ ;
wire \malu/Shift/_0439_ ;
wire \malu/Shift/_0440_ ;
wire \malu/Shift/_0441_ ;
wire \malu/Shift/_0442_ ;
wire \malu/Shift/_0443_ ;
wire \malu/Shift/_0444_ ;
wire \malu/Shift/_0445_ ;
wire \malu/Shift/_0446_ ;
wire \malu/Shift/_0447_ ;
wire \malu/Shift/_0448_ ;
wire \malu/Shift/_0449_ ;
wire \malu/Shift/_0450_ ;
wire \malu/Shift/_0451_ ;
wire \malu/Shift/_0452_ ;
wire \malu/Shift/_0453_ ;
wire \malu/Shift/_0454_ ;
wire \malu/Shift/_0455_ ;
wire \malu/Shift/_0456_ ;
wire \malu/Shift/_0457_ ;
wire \malu/Shift/_0458_ ;
wire \malu/Shift/_0459_ ;
wire \malu/Shift/_0460_ ;
wire \malu/Shift/_0461_ ;
wire \malu/Shift/_0462_ ;
wire \malu/Shift/_0463_ ;
wire \malu/Shift/_0464_ ;
wire \malu/Shift/_0465_ ;
wire \malu/Shift/_0466_ ;
wire \malu/Shift/_0467_ ;
wire \malu/Shift/_0468_ ;
wire \malu/Shift/_0469_ ;
wire \malu/Shift/_0470_ ;
wire \malu/Shift/_0471_ ;
wire \malu/Shift/_0472_ ;
wire \malu/Shift/_0473_ ;
wire \malu/Shift/_0474_ ;
wire \malu/Shift/_0475_ ;
wire \malu/Shift/_0476_ ;
wire \malu/Shift/_0477_ ;
wire \malu/Shift/_0478_ ;
wire \malu/Shift/_0479_ ;
wire \malu/Shift/_0480_ ;
wire \malu/Shift/_0481_ ;
wire \malu/Shift/_0482_ ;
wire \malu/Shift/_0483_ ;
wire \malu/Shift/_0484_ ;
wire \malu/Shift/_0485_ ;
wire \malu/Shift/_0486_ ;
wire \malu/Shift/_0487_ ;
wire \malu/Shift/_0488_ ;
wire \malu/Shift/_0489_ ;
wire \malu/Shift/_0490_ ;
wire \malu/Shift/_0491_ ;
wire \malu/Shift/_0492_ ;
wire \malu/Shift/_0493_ ;
wire \malu/Shift/_0494_ ;
wire \malu/Shift/_0495_ ;
wire \malu/Shift/_0496_ ;
wire \malu/Shift/_0497_ ;
wire \malu/Shift/_0498_ ;
wire \malu/Shift/_0499_ ;
wire \malu/Shift/_0500_ ;
wire \malu/Shift/_0501_ ;
wire \malu/Shift/_0502_ ;
wire \malu/Shift/_0503_ ;
wire \malu/Shift/_0504_ ;
wire \malu/Shift/_0505_ ;
wire \malu/Shift/_0506_ ;
wire \malu/Shift/_0507_ ;
wire \malu/Shift/_0508_ ;
wire \malu/Shift/_0509_ ;
wire \malu/Shift/_0510_ ;
wire \malu/Shift/_0511_ ;
wire \malu/Shift/_0512_ ;
wire \malu/Shift/_0513_ ;
wire \malu/Shift/_0514_ ;
wire \malu/Shift/_0515_ ;
wire \malu/Shift/_0516_ ;
wire \malu/Shift/_0517_ ;
wire \malu/Shift/_0518_ ;
wire \malu/Shift/_0519_ ;
wire \malu/Shift/_0520_ ;
wire \malu/Shift/_0521_ ;
wire \malu/Shift/_0522_ ;
wire \malu/Shift/_0523_ ;
wire \malu/Shift/_0524_ ;
wire \malu/Shift/_0525_ ;
wire \malu/Shift/_0526_ ;
wire \malu/Shift/_0527_ ;
wire \malu/Shift/_0528_ ;
wire \malu/Shift/_0529_ ;
wire \malu/Shift/_0530_ ;
wire \malu/Shift/_0531_ ;
wire \malu/Shift/_0532_ ;
wire \malu/Shift/_0533_ ;
wire \malu/Shift/_0534_ ;
wire \malu/Shift/_0535_ ;
wire \malu/Shift/_0536_ ;
wire \malu/Shift/_0537_ ;
wire \malu/Shift/_0538_ ;
wire \malu/Shift/_0539_ ;
wire \malu/Shift/_0540_ ;
wire \malu/Shift/_0541_ ;
wire \malu/Shift/_0542_ ;
wire \malu/Shift/_0543_ ;
wire \malu/Shift/_0544_ ;
wire \malu/Shift/_0545_ ;
wire \malu/Shift/_0546_ ;
wire \malu/Shift/_0547_ ;
wire \malu/Shift/_0548_ ;
wire \malu/Shift/_0549_ ;
wire \malu/Shift/_0550_ ;
wire \malu/Shift/_0551_ ;
wire \malu/Shift/_0552_ ;
wire \malu/Shift/_0553_ ;
wire \malu/Shift/_0554_ ;
wire \malu/Shift/_0555_ ;
wire \malu/Shift/_0556_ ;
wire \malu/Shift/_0557_ ;
wire \malu/Shift/_0558_ ;
wire \malu/Shift/_0559_ ;
wire \malu/Shift/_0560_ ;
wire \malu/Shift/_0561_ ;
wire \malu/Shift/_0562_ ;
wire \malu/Shift/_0563_ ;
wire \malu/Shift/_0564_ ;
wire \malu/Shift/_0565_ ;
wire \malu/Shift/_0566_ ;
wire \malu/Shift/_0567_ ;
wire \malu/Shift/_0568_ ;
wire \malu/Shift/_0569_ ;
wire \malu/Shift/_0570_ ;
wire \malu/Shift/_0571_ ;
wire \malu/Shift/_0572_ ;
wire \malu/Shift/_0573_ ;
wire \malu/Shift/_0574_ ;
wire \malu/Shift/_0575_ ;
wire \malu/Shift/_0576_ ;
wire \malu/Shift/_0577_ ;
wire \malu/Shift/_0578_ ;
wire \malu/Shift/_0579_ ;
wire \malu/Shift/_0580_ ;
wire \malu/Shift/_0581_ ;
wire \malu/Shift/_0582_ ;
wire \malu/Shift/_0583_ ;
wire \malu/Shift/_0584_ ;
wire \malu/Shift/_0585_ ;
wire \malu/Shift/_0586_ ;
wire \malu/Shift/_0587_ ;
wire \malu/Shift/_0588_ ;
wire \malu/Shift/_0589_ ;
wire \malu/Shift/_0590_ ;
wire \malu/Shift/_0591_ ;
wire \malu/Shift/_0592_ ;
wire \malu/Shift/_0593_ ;
wire \malu/Shift/_0594_ ;
wire \malu/Shift/_0595_ ;
wire \malu/Shift/_0596_ ;
wire \malu/Shift/_0597_ ;
wire \malu/Shift/_0598_ ;
wire \malu/Shift/_0599_ ;
wire \malu/Shift/_0600_ ;
wire \malu/Shift/_0601_ ;
wire \malu/Shift/_0602_ ;
wire \malu/Shift/_0603_ ;
wire \malu/Shift/_0604_ ;
wire \malu/Shift/_0605_ ;
wire \malu/Shift/_0606_ ;
wire \malu/Shift/_0607_ ;
wire \malu/Shift/_0608_ ;
wire \malu/Shift/_0609_ ;
wire \malu/Shift/_0610_ ;
wire \malu/Shift/_0611_ ;
wire \malu/Shift/_0612_ ;
wire \malu/Shift/_0613_ ;
wire \malu/Shift/_0614_ ;
wire \malu/Shift/_0615_ ;
wire \malu/Shift/_0616_ ;
wire \malu/Shift/_0617_ ;
wire \malu/Shift/_0618_ ;
wire \malu/Shift/_0619_ ;
wire \malu/Shift/_0620_ ;
wire \malu/Shift/_0621_ ;
wire \malu/Shift/_0622_ ;
wire \malu/Shift/_0623_ ;
wire \malu/Shift/_0624_ ;
wire \malu/Shift/_0625_ ;
wire \malu/Shift/_0626_ ;
wire \malu/Shift/_0627_ ;
wire \malu/Shift/_0628_ ;
wire \malu/Shift/_0629_ ;
wire \malu/Shift/_0630_ ;
wire \malu/Shift/_0631_ ;
wire \malu/Shift/_0632_ ;
wire \malu/Shift/_0633_ ;
wire \malu/Shift/_0634_ ;
wire \malu/Shift/_0635_ ;
wire \malu/Shift/_0636_ ;
wire \malu/Shift/_0637_ ;
wire \malu/Shift/_0638_ ;
wire \malu/Shift/_0639_ ;
wire \malu/Shift/_0640_ ;
wire \malu/Shift/_0641_ ;
wire \malu/Shift/_0642_ ;
wire \malu/Shift/_0643_ ;
wire \malu/Shift/_0644_ ;
wire \malu/Shift/_0645_ ;
wire \malu/Shift/_0646_ ;
wire \malu/Shift/_0647_ ;
wire \malu/Shift/_0648_ ;
wire \malu/Shift/_0649_ ;
wire \malu/Shift/_0650_ ;
wire \malu/Shift/_0651_ ;
wire \malu/Shift/_0652_ ;
wire \malu/Shift/_0653_ ;
wire \malu/Shift/_0654_ ;
wire \malu/Shift/_0655_ ;
wire \malu/Shift/_0656_ ;
wire \malu/Shift/_0657_ ;
wire \malu/Shift/_0658_ ;
wire \malu/Shift/_0659_ ;
wire \malu/Shift/_0660_ ;
wire \malu/Shift/_0661_ ;
wire \malu/Shift/_0662_ ;
wire \malu/Shift/_0663_ ;
wire \malu/Shift/_0664_ ;
wire \malu/Shift/_0665_ ;
wire \malu/Shift/_0666_ ;
wire \malu/Shift/_0667_ ;
wire \malu/Shift/_0668_ ;
wire \malu/Shift/_0669_ ;
wire \malu/Shift/_0670_ ;
wire \malu/Shift/_0671_ ;
wire \malu/Shift/_0672_ ;
wire \malu/Shift/_0673_ ;
wire \malu/Shift/_0674_ ;
wire \malu/Shift/_0675_ ;
wire \malu/Shift/_0676_ ;
wire \malu/Shift/_0677_ ;
wire \malu/Shift/_0678_ ;
wire \malu/Shift/_0679_ ;
wire \malu/Shift/_0680_ ;
wire \malu/Shift/_0681_ ;
wire \malu/Shift/_0682_ ;
wire \malu/Shift/_0683_ ;
wire \malu/Shift/_0684_ ;
wire \malu/Shift/_0685_ ;
wire \malu/Shift/_0686_ ;
wire \malu/Shift/_0687_ ;
wire \malu/Shift/_0688_ ;
wire \malu/Shift/_0689_ ;
wire \malu/Shift/_0690_ ;
wire \malu/Shift/_0691_ ;
wire \malu/Shift/_0692_ ;
wire \malu/Shift/_0693_ ;
wire \malu/Shift/_0694_ ;
wire \malu/Shift/_0695_ ;
wire \malu/Shift/_0696_ ;
wire \malu/Shift/_0697_ ;
wire \malu/Shift/_0698_ ;
wire \malu/Shift/_0699_ ;
wire \malu/Shift/_0700_ ;
wire \malu/Shift/_0701_ ;
wire \malu/Shift/_0702_ ;
wire \malu/Shift/_0703_ ;
wire \malu/Shift/_0704_ ;
wire \malu/Shift/_0705_ ;
wire \malu/Shift/_0706_ ;
wire \malu/Shift/_0707_ ;
wire \malu/Shift/_0708_ ;
wire \malu/Shift/_0709_ ;
wire \malu/Shift/_0710_ ;
wire \malu/Shift/_0711_ ;
wire \malu/Shift/_0712_ ;
wire \malu/Shift/_0713_ ;
wire \malu/Shift/_0714_ ;
wire \malu/Shift/_0715_ ;
wire \malu/Shift/_0716_ ;
wire \malu/Shift/_0717_ ;
wire \malu/Shift/_0718_ ;
wire \malu/Shift/_0719_ ;
wire \malu/Shift/_0720_ ;
wire \malu/Shift/_0721_ ;
wire \malu/Shift/_0722_ ;
wire \malu/Shift/_0723_ ;
wire \malu/Shift/_0724_ ;
wire \malu/Shift/_0725_ ;
wire \malu/Shift/_0726_ ;
wire \malu/Shift/_0727_ ;
wire \malu/Shift/_0728_ ;
wire \malu/Shift/_0729_ ;
wire \malu/Shift/_0730_ ;
wire \malu/Shift/_0731_ ;
wire \malu/Shift/_0732_ ;
wire \malu/Shift/_0733_ ;
wire \malu/Shift/_0734_ ;
wire \malu/Shift/_0735_ ;
wire \malu/Shift/_0736_ ;
wire \malu/Shift/_0737_ ;
wire \malu/Shift/_0738_ ;
wire \malu/Shift/_0739_ ;
wire \malu/Shift/_0740_ ;
wire \malu/Shift/_0741_ ;
wire \malu/Shift/_0742_ ;
wire \malu/Shift/_0743_ ;
wire \malu/Shift/_0744_ ;
wire \malu/Shift/_0745_ ;
wire \malu/Shift/_0746_ ;
wire \malu/Shift/_0747_ ;
wire \malu/Shift/_0748_ ;
wire \malu/Shift/_0749_ ;
wire \malu/Shift/_0750_ ;
wire \malu/Shift/_0751_ ;
wire \malu/Shift/_0752_ ;
wire \marbiter/_0000_ ;
wire \marbiter/_0001_ ;
wire \marbiter/_0002_ ;
wire \marbiter/_0003_ ;
wire \marbiter/_0004_ ;
wire \marbiter/_0005_ ;
wire \marbiter/_0006_ ;
wire \marbiter/_0007_ ;
wire \marbiter/_0008_ ;
wire \marbiter/_0009_ ;
wire \marbiter/_0010_ ;
wire \marbiter/_0011_ ;
wire \marbiter/_0012_ ;
wire \marbiter/_0013_ ;
wire \marbiter/_0014_ ;
wire \marbiter/_0015_ ;
wire \marbiter/_0016_ ;
wire \marbiter/_0017_ ;
wire \marbiter/_0018_ ;
wire \marbiter/_0019_ ;
wire \marbiter/_0020_ ;
wire \marbiter/_0021_ ;
wire \marbiter/_0022_ ;
wire \marbiter/_0023_ ;
wire \marbiter/_0024_ ;
wire \marbiter/_0025_ ;
wire \marbiter/_0026_ ;
wire \marbiter/_0027_ ;
wire \marbiter/_0028_ ;
wire \marbiter/_0029_ ;
wire \marbiter/_0030_ ;
wire \marbiter/_0031_ ;
wire \marbiter/_0032_ ;
wire \marbiter/_0033_ ;
wire \marbiter/_0034_ ;
wire \marbiter/_0035_ ;
wire \marbiter/_0036_ ;
wire \marbiter/_0037_ ;
wire \marbiter/_0038_ ;
wire \marbiter/_0039_ ;
wire \marbiter/_0040_ ;
wire \marbiter/_0041_ ;
wire \marbiter/_0042_ ;
wire \marbiter/_0043_ ;
wire \marbiter/_0044_ ;
wire \marbiter/_0045_ ;
wire \marbiter/_0046_ ;
wire \marbiter/_0047_ ;
wire \marbiter/_0048_ ;
wire \marbiter/_0049_ ;
wire \marbiter/_0050_ ;
wire \marbiter/_0051_ ;
wire \marbiter/_0052_ ;
wire \marbiter/_0053_ ;
wire \marbiter/_0054_ ;
wire \marbiter/_0055_ ;
wire \marbiter/_0056_ ;
wire \marbiter/_0057_ ;
wire \marbiter/_0058_ ;
wire \marbiter/_0059_ ;
wire \marbiter/_0060_ ;
wire \marbiter/_0061_ ;
wire \marbiter/_0062_ ;
wire \marbiter/_0063_ ;
wire \marbiter/_0064_ ;
wire \marbiter/_0065_ ;
wire \marbiter/_0066_ ;
wire \marbiter/_0067_ ;
wire \marbiter/_0068_ ;
wire \marbiter/_0069_ ;
wire \marbiter/_0070_ ;
wire \marbiter/_0071_ ;
wire \marbiter/_0072_ ;
wire \marbiter/_0073_ ;
wire \marbiter/_0074_ ;
wire \marbiter/_0075_ ;
wire \marbiter/_0076_ ;
wire \marbiter/_0077_ ;
wire \marbiter/_0078_ ;
wire \marbiter/_0079_ ;
wire \marbiter/_0080_ ;
wire \marbiter/_0081_ ;
wire \marbiter/_0082_ ;
wire \marbiter/_0083_ ;
wire \marbiter/_0084_ ;
wire \marbiter/_0085_ ;
wire \marbiter/_0086_ ;
wire \marbiter/_0087_ ;
wire \marbiter/_0088_ ;
wire \marbiter/_0089_ ;
wire \marbiter/_0090_ ;
wire \marbiter/_0091_ ;
wire \marbiter/_0092_ ;
wire \marbiter/_0093_ ;
wire \marbiter/_0094_ ;
wire \marbiter/_0095_ ;
wire \marbiter/_0096_ ;
wire \marbiter/_0097_ ;
wire \marbiter/_0098_ ;
wire \marbiter/_0099_ ;
wire \marbiter/_0100_ ;
wire \marbiter/_0101_ ;
wire \marbiter/_0102_ ;
wire \marbiter/_0103_ ;
wire \marbiter/_0104_ ;
wire \marbiter/_0105_ ;
wire \marbiter/_0106_ ;
wire \marbiter/_0107_ ;
wire \marbiter/_0108_ ;
wire \marbiter/_0109_ ;
wire \marbiter/_0110_ ;
wire \marbiter/_0111_ ;
wire \marbiter/_0112_ ;
wire \marbiter/_0113_ ;
wire \marbiter/_0114_ ;
wire \marbiter/_0115_ ;
wire \marbiter/_0116_ ;
wire \marbiter/_0117_ ;
wire \marbiter/_0118_ ;
wire \marbiter/_0119_ ;
wire \marbiter/_0120_ ;
wire \marbiter/_0121_ ;
wire \marbiter/_0122_ ;
wire \marbiter/_0123_ ;
wire \marbiter/_0124_ ;
wire \marbiter/_0125_ ;
wire \marbiter/_0126_ ;
wire \marbiter/_0127_ ;
wire \marbiter/_0128_ ;
wire \marbiter/_0129_ ;
wire \marbiter/_0130_ ;
wire \marbiter/_0131_ ;
wire \marbiter/_0132_ ;
wire \marbiter/_0133_ ;
wire \marbiter/_0134_ ;
wire \marbiter/_0135_ ;
wire \marbiter/_0136_ ;
wire \marbiter/_0137_ ;
wire \marbiter/_0138_ ;
wire \marbiter/_0139_ ;
wire \marbiter/_0140_ ;
wire \marbiter/_0141_ ;
wire \marbiter/_0142_ ;
wire \marbiter/_0143_ ;
wire \marbiter/_0144_ ;
wire \marbiter/_0145_ ;
wire \marbiter/_0146_ ;
wire \marbiter/_0147_ ;
wire \marbiter/_0148_ ;
wire \marbiter/_0149_ ;
wire \marbiter/_0150_ ;
wire \marbiter/_0151_ ;
wire \marbiter/_0152_ ;
wire \marbiter/_0153_ ;
wire \marbiter/_0154_ ;
wire \marbiter/_0155_ ;
wire \marbiter/_0156_ ;
wire \marbiter/_0157_ ;
wire \marbiter/_0158_ ;
wire \marbiter/_0159_ ;
wire \marbiter/_0160_ ;
wire \marbiter/_0161_ ;
wire \marbiter/_0162_ ;
wire \marbiter/_0163_ ;
wire \marbiter/_0164_ ;
wire \marbiter/_0165_ ;
wire \marbiter/_0166_ ;
wire \marbiter/_0167_ ;
wire \marbiter/_0168_ ;
wire \marbiter/_0169_ ;
wire \marbiter/_0170_ ;
wire \marbiter/_0171_ ;
wire \marbiter/_0172_ ;
wire \marbiter/_0173_ ;
wire \marbiter/_0174_ ;
wire \marbiter/_0175_ ;
wire \marbiter/_0176_ ;
wire \marbiter/_0177_ ;
wire \marbiter/_0178_ ;
wire \marbiter/_0179_ ;
wire \marbiter/_0180_ ;
wire \marbiter/_0181_ ;
wire \marbiter/_0182_ ;
wire \marbiter/_0183_ ;
wire \marbiter/_0184_ ;
wire \marbiter/_0185_ ;
wire \marbiter/_0186_ ;
wire \marbiter/_0187_ ;
wire \marbiter/_0188_ ;
wire \marbiter/_0189_ ;
wire \marbiter/_0190_ ;
wire \marbiter/_0191_ ;
wire \marbiter/_0192_ ;
wire \marbiter/_0193_ ;
wire \marbiter/_0194_ ;
wire \marbiter/_0195_ ;
wire \marbiter/_0196_ ;
wire \marbiter/_0197_ ;
wire \marbiter/_0198_ ;
wire \marbiter/_0199_ ;
wire \marbiter/_0200_ ;
wire \marbiter/_0201_ ;
wire \marbiter/_0202_ ;
wire \marbiter/_0203_ ;
wire \marbiter/_0204_ ;
wire \marbiter/_0205_ ;
wire \marbiter/_0206_ ;
wire \marbiter/_0207_ ;
wire \marbiter/_0208_ ;
wire \marbiter/_0209_ ;
wire \marbiter/_0210_ ;
wire \marbiter/_0211_ ;
wire \marbiter/_0212_ ;
wire \marbiter/_0213_ ;
wire \marbiter/_0214_ ;
wire \marbiter/_0215_ ;
wire \marbiter/_0216_ ;
wire \marbiter/_0217_ ;
wire \marbiter/_0218_ ;
wire \marbiter/_0219_ ;
wire \marbiter/_0220_ ;
wire \marbiter/_0221_ ;
wire \marbiter/_0222_ ;
wire \marbiter/_0223_ ;
wire \marbiter/_0224_ ;
wire \marbiter/_0225_ ;
wire \marbiter/_0226_ ;
wire \marbiter/_0227_ ;
wire \marbiter/_0228_ ;
wire \marbiter/_0229_ ;
wire \marbiter/_0230_ ;
wire \marbiter/_0231_ ;
wire \marbiter/_0232_ ;
wire \marbiter/_0233_ ;
wire \marbiter/_0234_ ;
wire \marbiter/_0235_ ;
wire \marbiter/_0236_ ;
wire \marbiter/_0237_ ;
wire \marbiter/_0238_ ;
wire \marbiter/_0239_ ;
wire \marbiter/_0240_ ;
wire \marbiter/_0241_ ;
wire \marbiter/_0242_ ;
wire \marbiter/_0243_ ;
wire \marbiter/_0244_ ;
wire \marbiter/_0245_ ;
wire \marbiter/_0246_ ;
wire \marbiter/_0247_ ;
wire \marbiter/_0248_ ;
wire \marbiter/_0249_ ;
wire \marbiter/_0250_ ;
wire \marbiter/_0251_ ;
wire \marbiter/_0252_ ;
wire \marbiter/_0253_ ;
wire \marbiter/_0254_ ;
wire \marbiter/_0255_ ;
wire \marbiter/_0256_ ;
wire \marbiter/_0257_ ;
wire \marbiter/_0258_ ;
wire \marbiter/_0259_ ;
wire \marbiter/_0260_ ;
wire \marbiter/_0261_ ;
wire \marbiter/_0262_ ;
wire \marbiter/_0263_ ;
wire \marbiter/_0264_ ;
wire \marbiter/_0265_ ;
wire \marbiter/_0266_ ;
wire \marbiter/_0267_ ;
wire \marbiter/_0268_ ;
wire \marbiter/_0269_ ;
wire \marbiter/_0270_ ;
wire \marbiter/_0271_ ;
wire \marbiter/_0272_ ;
wire \marbiter/_0273_ ;
wire \marbiter/_0274_ ;
wire \marbiter/_0275_ ;
wire \marbiter/_0276_ ;
wire \marbiter/_0277_ ;
wire \marbiter/_0278_ ;
wire \marbiter/_0279_ ;
wire \marbiter/_0280_ ;
wire \marbiter/_0281_ ;
wire \marbiter/_0282_ ;
wire \marbiter/_0283_ ;
wire \marbiter/_0284_ ;
wire \marbiter/_0285_ ;
wire \marbiter/_0286_ ;
wire \marbiter/_0287_ ;
wire \marbiter/_0288_ ;
wire \marbiter/_0289_ ;
wire \marbiter/_0290_ ;
wire \marbiter/_0291_ ;
wire \marbiter/_0292_ ;
wire \marbiter/_0293_ ;
wire \marbiter/_0294_ ;
wire \marbiter/_0295_ ;
wire \marbiter/_0296_ ;
wire \marbiter/_0297_ ;
wire \marbiter/_0298_ ;
wire \marbiter/_0299_ ;
wire \marbiter/_0300_ ;
wire \marbiter/_0301_ ;
wire \marbiter/_0302_ ;
wire \marbiter/_0303_ ;
wire \marbiter/_0304_ ;
wire \marbiter/_0305_ ;
wire \marbiter/_0306_ ;
wire \marbiter/_0307_ ;
wire \marbiter/_0308_ ;
wire \marbiter/_0309_ ;
wire \marbiter/_0310_ ;
wire \marbiter/_0311_ ;
wire \marbiter/_0312_ ;
wire \marbiter/_0313_ ;
wire \marbiter/_0314_ ;
wire \marbiter/_0315_ ;
wire \marbiter/_0316_ ;
wire \marbiter/_0317_ ;
wire \marbiter/_0318_ ;
wire \marbiter/_0319_ ;
wire \marbiter/_0320_ ;
wire \marbiter/_0321_ ;
wire \marbiter/_0322_ ;
wire \marbiter/_0323_ ;
wire \marbiter/_0324_ ;
wire \marbiter/_0325_ ;
wire \marbiter/_0326_ ;
wire \marbiter/_0327_ ;
wire \marbiter/_0328_ ;
wire \marbiter/_0329_ ;
wire \marbiter/_0330_ ;
wire \marbiter/_0331_ ;
wire \marbiter/_0332_ ;
wire \marbiter/_0333_ ;
wire \marbiter/_0334_ ;
wire \marbiter/_0335_ ;
wire \marbiter/_0336_ ;
wire \marbiter/_0337_ ;
wire \marbiter/_0338_ ;
wire \marbiter/_0339_ ;
wire \marbiter/_0340_ ;
wire \marbiter/_0341_ ;
wire \marbiter/_0342_ ;
wire \marbiter/_0343_ ;
wire \marbiter/_0344_ ;
wire \marbiter/_0345_ ;
wire \marbiter/_0346_ ;
wire \marbiter/_0347_ ;
wire \marbiter/_0348_ ;
wire \marbiter/_0349_ ;
wire \marbiter/_0350_ ;
wire \marbiter/_0351_ ;
wire \marbiter/_0352_ ;
wire \marbiter/_0353_ ;
wire \marbiter/_0354_ ;
wire \marbiter/_0355_ ;
wire \marbiter/_0356_ ;
wire \marbiter/_0357_ ;
wire \marbiter/_0358_ ;
wire \marbiter/_0359_ ;
wire \marbiter/_0360_ ;
wire \marbiter/_0361_ ;
wire \marbiter/_0362_ ;
wire \marbiter/_0363_ ;
wire \marbiter/_0364_ ;
wire \marbiter/_0365_ ;
wire \marbiter/_0366_ ;
wire \marbiter/_0367_ ;
wire \marbiter/_0368_ ;
wire \marbiter/_0369_ ;
wire \marbiter/_0370_ ;
wire \marbiter/_0371_ ;
wire \marbiter/_0372_ ;
wire \marbiter/_0373_ ;
wire \marbiter/_0374_ ;
wire \marbiter/_0375_ ;
wire \marbiter/_0376_ ;
wire \marbiter/_0377_ ;
wire \marbiter/_0378_ ;
wire \marbiter/_0379_ ;
wire \marbiter/_0380_ ;
wire \marbiter/_0381_ ;
wire \marbiter/_0382_ ;
wire \marbiter/_0383_ ;
wire \marbiter/_0384_ ;
wire \marbiter/_0385_ ;
wire \marbiter/_0386_ ;
wire \marbiter/_0387_ ;
wire \marbiter/_0388_ ;
wire \marbiter/_0389_ ;
wire \marbiter/_0390_ ;
wire \marbiter/_0391_ ;
wire \marbiter/_0392_ ;
wire \marbiter/_0393_ ;
wire \marbiter/_0394_ ;
wire \marbiter/_0395_ ;
wire \marbiter/_0396_ ;
wire \marbiter/_0397_ ;
wire \marbiter/_0398_ ;
wire \marbiter/_0399_ ;
wire \marbiter/_0400_ ;
wire \marbiter/_0401_ ;
wire \marbiter/_0402_ ;
wire \marbiter/_0403_ ;
wire \marbiter/_0404_ ;
wire \marbiter/_0405_ ;
wire \marbiter/_0406_ ;
wire \marbiter/_0407_ ;
wire \marbiter/_0408_ ;
wire \marbiter/_0409_ ;
wire \marbiter/_0410_ ;
wire \marbiter/_0411_ ;
wire \marbiter/_0412_ ;
wire \marbiter/_0413_ ;
wire \marbiter/_0414_ ;
wire \marbiter/_0415_ ;
wire \marbiter/_0416_ ;
wire \marbiter/_0417_ ;
wire \marbiter/_0418_ ;
wire \marbiter/_0419_ ;
wire \marbiter/_0420_ ;
wire \marbiter/_0421_ ;
wire \marbiter/_0422_ ;
wire \marbiter/_0423_ ;
wire \marbiter/_0424_ ;
wire \marbiter/_0425_ ;
wire \marbiter/_0426_ ;
wire \marbiter/_0427_ ;
wire \marbiter/_0428_ ;
wire \marbiter/_0429_ ;
wire \marbiter/_0430_ ;
wire \marbiter/_0431_ ;
wire \marbiter/_0432_ ;
wire \marbiter/_0433_ ;
wire \marbiter/_0434_ ;
wire \marbiter/_0435_ ;
wire \marbiter/_0436_ ;
wire \marbiter/_0437_ ;
wire \marbiter/_0438_ ;
wire \marbiter/_0439_ ;
wire \marbiter/_0440_ ;
wire \marbiter/_0441_ ;
wire \marbiter/_0442_ ;
wire \marbiter/_0443_ ;
wire \marbiter/_0444_ ;
wire \marbiter/_0445_ ;
wire \marbiter/_0446_ ;
wire \marbiter/_0447_ ;
wire \marbiter/_0448_ ;
wire \marbiter/_0449_ ;
wire \marbiter/_0450_ ;
wire \marbiter/_0451_ ;
wire \marbiter/_0452_ ;
wire \marbiter/_0453_ ;
wire \marbiter/_0454_ ;
wire \marbiter/_0455_ ;
wire \marbiter/_0456_ ;
wire \marbiter/_0457_ ;
wire \marbiter/_0458_ ;
wire \marbiter/_0459_ ;
wire \marbiter/_0460_ ;
wire \marbiter/_0461_ ;
wire \marbiter/_0462_ ;
wire \marbiter/_0463_ ;
wire \marbiter/_0464_ ;
wire \marbiter/_0465_ ;
wire \marbiter/_0466_ ;
wire \marbiter/_0467_ ;
wire \marbiter/_0468_ ;
wire \marbiter/_0469_ ;
wire \marbiter/_0470_ ;
wire \marbiter/_0471_ ;
wire \marbiter/_0472_ ;
wire \marbiter/_0473_ ;
wire \marbiter/_0474_ ;
wire \marbiter/_0475_ ;
wire \marbiter/_0476_ ;
wire \marbiter/_0477_ ;
wire \marbiter/_0478_ ;
wire \marbiter/_0479_ ;
wire \marbiter/_0480_ ;
wire \marbiter/_0481_ ;
wire \marbiter/_0482_ ;
wire \marbiter/_0483_ ;
wire \marbiter/_0484_ ;
wire \marbiter/_0485_ ;
wire \marbiter/_0486_ ;
wire \marbiter/_0487_ ;
wire \marbiter/_0488_ ;
wire \marbiter/_0489_ ;
wire \marbiter/_0490_ ;
wire \marbiter/_0491_ ;
wire \marbiter/_0492_ ;
wire \marbiter/_0493_ ;
wire \marbiter/_0494_ ;
wire \marbiter/_0495_ ;
wire \marbiter/_0496_ ;
wire \marbiter/_0497_ ;
wire \marbiter/_0498_ ;
wire \marbiter/_0499_ ;
wire \marbiter/_0500_ ;
wire \marbiter/_0501_ ;
wire \marbiter/_0502_ ;
wire \marbiter/_0503_ ;
wire \marbiter/_0504_ ;
wire \marbiter/_0505_ ;
wire \marbiter/_0506_ ;
wire \marbiter/_0507_ ;
wire \marbiter/_0508_ ;
wire \marbiter/_0509_ ;
wire \marbiter/_0510_ ;
wire \marbiter/_0511_ ;
wire \marbiter/_0512_ ;
wire \marbiter/_0513_ ;
wire \marbiter/_0514_ ;
wire \marbiter/_0515_ ;
wire \marbiter/_0516_ ;
wire \marbiter/_0517_ ;
wire \marbiter/_0518_ ;
wire \marbiter/_0519_ ;
wire \marbiter/_0520_ ;
wire \marbiter/_0521_ ;
wire \marbiter/_0522_ ;
wire \marbiter/_0523_ ;
wire \marbiter/_0524_ ;
wire \marbiter/_0525_ ;
wire \marbiter/_0526_ ;
wire \marbiter/_0527_ ;
wire \marbiter/_0528_ ;
wire \marbiter/_0529_ ;
wire \marbiter/_0530_ ;
wire \marbiter/_0531_ ;
wire \marbiter/_0532_ ;
wire \marbiter/_0533_ ;
wire \marbiter/_0534_ ;
wire \marbiter/_0535_ ;
wire \marbiter/_0536_ ;
wire \marbiter/_0537_ ;
wire \marbiter/_0538_ ;
wire \marbiter/_0539_ ;
wire \marbiter/_0540_ ;
wire \marbiter/_0541_ ;
wire \marbiter/_0542_ ;
wire \marbiter/_0543_ ;
wire \marbiter/_0544_ ;
wire \marbiter/_0545_ ;
wire \marbiter/_0546_ ;
wire \marbiter/_0547_ ;
wire \marbiter/_0548_ ;
wire \marbiter/_0549_ ;
wire \marbiter/_0550_ ;
wire \marbiter/_0551_ ;
wire \marbiter/_0552_ ;
wire \marbiter/_0553_ ;
wire \marbiter/_0554_ ;
wire \marbiter/_0555_ ;
wire \marbiter/_0556_ ;
wire \marbiter/_0557_ ;
wire \marbiter/_0558_ ;
wire \marbiter/_0559_ ;
wire \marbiter/_0560_ ;
wire \marbiter/_0561_ ;
wire \marbiter/_0562_ ;
wire \marbiter/_0563_ ;
wire \marbiter/_0564_ ;
wire \marbiter/_0565_ ;
wire \marbiter/_0566_ ;
wire \marbiter/_0567_ ;
wire \marbiter/_0568_ ;
wire \marbiter/_0569_ ;
wire \marbiter/_0570_ ;
wire \marbiter/_0571_ ;
wire \marbiter/_0572_ ;
wire \marbiter/_0573_ ;
wire \marbiter/_0574_ ;
wire \marbiter/_0575_ ;
wire \marbiter/_0576_ ;
wire \marbiter/_0577_ ;
wire \marbiter/_0578_ ;
wire \marbiter/_0579_ ;
wire \marbiter/_0580_ ;
wire \marbiter/_0581_ ;
wire \marbiter/_0582_ ;
wire \marbiter/_0583_ ;
wire \marbiter/_0584_ ;
wire \marbiter/_0585_ ;
wire \marbiter/_0586_ ;
wire \marbiter/_0587_ ;
wire \marbiter/_0588_ ;
wire \marbiter/_0589_ ;
wire \marbiter/_0590_ ;
wire \marbiter/_0591_ ;
wire \marbiter/_0592_ ;
wire \marbiter/_0593_ ;
wire \marbiter/_0594_ ;
wire \marbiter/_0595_ ;
wire \marbiter/_0596_ ;
wire \marbiter/_0597_ ;
wire \marbiter/_0598_ ;
wire \marbiter/_0599_ ;
wire \marbiter/_0600_ ;
wire \marbiter/_0601_ ;
wire \marbiter/_0602_ ;
wire \marbiter/_0603_ ;
wire \marbiter/_0604_ ;
wire \marbiter/_0605_ ;
wire \marbiter/_0606_ ;
wire \marbiter/_0607_ ;
wire \marbiter/_0608_ ;
wire \marbiter/_0609_ ;
wire \marbiter/_0610_ ;
wire \marbiter/_0611_ ;
wire \marbiter/_0612_ ;
wire \marbiter/_0613_ ;
wire \marbiter/_0614_ ;
wire \marbiter/_0615_ ;
wire \marbiter/_0616_ ;
wire \marbiter/_0617_ ;
wire \marbiter/_0618_ ;
wire \marbiter/_0619_ ;
wire \marbiter/_0620_ ;
wire \marbiter/_0621_ ;
wire \marbiter/_0622_ ;
wire \marbiter/_0623_ ;
wire \marbiter/_0624_ ;
wire \marbiter/_0625_ ;
wire \marbiter/_0626_ ;
wire \marbiter/_0627_ ;
wire \marbiter/_0628_ ;
wire \marbiter/_0629_ ;
wire \marbiter/_0630_ ;
wire \marbiter/_0631_ ;
wire \marbiter/_0632_ ;
wire \marbiter/_0633_ ;
wire \marbiter/_0634_ ;
wire \marbiter/_0635_ ;
wire \marbiter/_0636_ ;
wire \marbiter/_0637_ ;
wire \marbiter/_0638_ ;
wire \marbiter/_0639_ ;
wire \marbiter/_0640_ ;
wire \marbiter/_0641_ ;
wire \marbiter/_0642_ ;
wire \marbiter/_0643_ ;
wire \marbiter/_0644_ ;
wire \marbiter/_0645_ ;
wire \marbiter/_0646_ ;
wire \marbiter/_0647_ ;
wire \marbiter/_0648_ ;
wire \marbiter/_0649_ ;
wire \marbiter/_0650_ ;
wire \marbiter/_0651_ ;
wire \marbiter/_0652_ ;
wire \marbiter/_0653_ ;
wire \marbiter/_0654_ ;
wire \marbiter/_0655_ ;
wire \marbiter/_0656_ ;
wire \marbiter/_0657_ ;
wire \marbiter/_0658_ ;
wire \marbiter/_0659_ ;
wire \marbiter/_0660_ ;
wire \marbiter/_0661_ ;
wire \marbiter/_0662_ ;
wire \marbiter/_0663_ ;
wire \marbiter/_0664_ ;
wire \marbiter/_0665_ ;
wire \marbiter/_0666_ ;
wire \marbiter/_0667_ ;
wire \marbiter/_0668_ ;
wire \marbiter/_0669_ ;
wire \marbiter/_0670_ ;
wire \marbiter/_0671_ ;
wire \marbiter/_0672_ ;
wire \marbiter/_0673_ ;
wire \marbiter/_0674_ ;
wire \marbiter/_0675_ ;
wire \marbiter/_0676_ ;
wire \marbiter/_0677_ ;
wire \marbiter/_0678_ ;
wire \marbiter/_0679_ ;
wire \marbiter/_0680_ ;
wire \marbiter/_0681_ ;
wire \marbiter/_0682_ ;
wire \marbiter/_0683_ ;
wire \marbiter/_0684_ ;
wire \marbiter/_0685_ ;
wire \marbiter/_0686_ ;
wire \marbiter/_0687_ ;
wire \marbiter/_0688_ ;
wire \marbiter/_0689_ ;
wire \marbiter/_0690_ ;
wire \marbiter/_0691_ ;
wire \marbiter/_0692_ ;
wire \marbiter/_0693_ ;
wire \marbiter/_0694_ ;
wire \marbiter/_0695_ ;
wire \marbiter/_0696_ ;
wire \marbiter/_0697_ ;
wire \marbiter/_0698_ ;
wire \marbiter/_0699_ ;
wire \marbiter/_0700_ ;
wire \marbiter/_0701_ ;
wire \marbiter/_0702_ ;
wire \marbiter/_0703_ ;
wire \marbiter/_0704_ ;
wire \marbiter/_0705_ ;
wire \marbiter/_0706_ ;
wire \marbiter/_0707_ ;
wire \marbiter/_0708_ ;
wire \marbiter/_0709_ ;
wire \marbiter/read_state[0] ;
wire \marbiter/read_state[1] ;
wire \marbiter/read_state[2] ;
wire \marbiter/write_state[0] ;
wire \marbiter/write_state[1] ;
wire \marbiter/write_state[2] ;
wire \mcsr/_0000_ ;
wire \mcsr/_0001_ ;
wire \mcsr/_0002_ ;
wire \mcsr/_0003_ ;
wire \mcsr/_0004_ ;
wire \mcsr/_0005_ ;
wire \mcsr/_0006_ ;
wire \mcsr/_0007_ ;
wire \mcsr/_0008_ ;
wire \mcsr/_0009_ ;
wire \mcsr/_0010_ ;
wire \mcsr/_0011_ ;
wire \mcsr/_0012_ ;
wire \mcsr/_0013_ ;
wire \mcsr/_0014_ ;
wire \mcsr/_0015_ ;
wire \mcsr/_0016_ ;
wire \mcsr/_0017_ ;
wire \mcsr/_0018_ ;
wire \mcsr/_0019_ ;
wire \mcsr/_0020_ ;
wire \mcsr/_0021_ ;
wire \mcsr/_0022_ ;
wire \mcsr/_0023_ ;
wire \mcsr/_0024_ ;
wire \mcsr/_0025_ ;
wire \mcsr/_0026_ ;
wire \mcsr/_0027_ ;
wire \mcsr/_0028_ ;
wire \mcsr/_0029_ ;
wire \mcsr/_0030_ ;
wire \mcsr/_0031_ ;
wire \mcsr/_0032_ ;
wire \mcsr/_0033_ ;
wire \mcsr/_0034_ ;
wire \mcsr/_0035_ ;
wire \mcsr/_0036_ ;
wire \mcsr/_0037_ ;
wire \mcsr/_0038_ ;
wire \mcsr/_0039_ ;
wire \mcsr/_0040_ ;
wire \mcsr/_0041_ ;
wire \mcsr/_0042_ ;
wire \mcsr/_0043_ ;
wire \mcsr/_0044_ ;
wire \mcsr/_0045_ ;
wire \mcsr/_0046_ ;
wire \mcsr/_0047_ ;
wire \mcsr/_0048_ ;
wire \mcsr/_0049_ ;
wire \mcsr/_0050_ ;
wire \mcsr/_0051_ ;
wire \mcsr/_0052_ ;
wire \mcsr/_0053_ ;
wire \mcsr/_0054_ ;
wire \mcsr/_0055_ ;
wire \mcsr/_0056_ ;
wire \mcsr/_0057_ ;
wire \mcsr/_0058_ ;
wire \mcsr/_0059_ ;
wire \mcsr/_0060_ ;
wire \mcsr/_0061_ ;
wire \mcsr/_0062_ ;
wire \mcsr/_0063_ ;
wire \mcsr/_0064_ ;
wire \mcsr/_0065_ ;
wire \mcsr/_0066_ ;
wire \mcsr/_0067_ ;
wire \mcsr/_0068_ ;
wire \mcsr/_0069_ ;
wire \mcsr/_0070_ ;
wire \mcsr/_0071_ ;
wire \mcsr/_0072_ ;
wire \mcsr/_0073_ ;
wire \mcsr/_0074_ ;
wire \mcsr/_0075_ ;
wire \mcsr/_0076_ ;
wire \mcsr/_0077_ ;
wire \mcsr/_0078_ ;
wire \mcsr/_0079_ ;
wire \mcsr/_0080_ ;
wire \mcsr/_0081_ ;
wire \mcsr/_0082_ ;
wire \mcsr/_0083_ ;
wire \mcsr/_0084_ ;
wire \mcsr/_0085_ ;
wire \mcsr/_0086_ ;
wire \mcsr/_0087_ ;
wire \mcsr/_0088_ ;
wire \mcsr/_0089_ ;
wire \mcsr/_0090_ ;
wire \mcsr/_0091_ ;
wire \mcsr/_0092_ ;
wire \mcsr/_0093_ ;
wire \mcsr/_0094_ ;
wire \mcsr/_0095_ ;
wire \mcsr/_0096_ ;
wire \mcsr/_0097_ ;
wire \mcsr/_0098_ ;
wire \mcsr/_0099_ ;
wire \mcsr/_0100_ ;
wire \mcsr/_0101_ ;
wire \mcsr/_0102_ ;
wire \mcsr/_0103_ ;
wire \mcsr/_0104_ ;
wire \mcsr/_0105_ ;
wire \mcsr/_0106_ ;
wire \mcsr/_0107_ ;
wire \mcsr/_0108_ ;
wire \mcsr/_0109_ ;
wire \mcsr/_0110_ ;
wire \mcsr/_0111_ ;
wire \mcsr/_0112_ ;
wire \mcsr/_0113_ ;
wire \mcsr/_0114_ ;
wire \mcsr/_0115_ ;
wire \mcsr/_0116_ ;
wire \mcsr/_0117_ ;
wire \mcsr/_0118_ ;
wire \mcsr/_0119_ ;
wire \mcsr/_0120_ ;
wire \mcsr/_0121_ ;
wire \mcsr/_0122_ ;
wire \mcsr/_0123_ ;
wire \mcsr/_0124_ ;
wire \mcsr/_0125_ ;
wire \mcsr/_0126_ ;
wire \mcsr/_0127_ ;
wire \mcsr/_0128_ ;
wire \mcsr/_0129_ ;
wire \mcsr/_0130_ ;
wire \mcsr/_0131_ ;
wire \mcsr/_0132_ ;
wire \mcsr/_0133_ ;
wire \mcsr/_0134_ ;
wire \mcsr/_0135_ ;
wire \mcsr/_0136_ ;
wire \mcsr/_0137_ ;
wire \mcsr/_0138_ ;
wire \mcsr/_0139_ ;
wire \mcsr/_0140_ ;
wire \mcsr/_0141_ ;
wire \mcsr/_0142_ ;
wire \mcsr/_0143_ ;
wire \mcsr/_0144_ ;
wire \mcsr/_0145_ ;
wire \mcsr/_0146_ ;
wire \mcsr/_0147_ ;
wire \mcsr/_0148_ ;
wire \mcsr/_0149_ ;
wire \mcsr/_0150_ ;
wire \mcsr/_0151_ ;
wire \mcsr/_0152_ ;
wire \mcsr/_0153_ ;
wire \mcsr/_0154_ ;
wire \mcsr/_0155_ ;
wire \mcsr/_0156_ ;
wire \mcsr/_0157_ ;
wire \mcsr/_0158_ ;
wire \mcsr/_0159_ ;
wire \mcsr/_0160_ ;
wire \mcsr/_0161_ ;
wire \mcsr/_0162_ ;
wire \mcsr/_0163_ ;
wire \mcsr/_0164_ ;
wire \mcsr/_0165_ ;
wire \mcsr/_0166_ ;
wire \mcsr/_0167_ ;
wire \mcsr/_0168_ ;
wire \mcsr/_0169_ ;
wire \mcsr/_0170_ ;
wire \mcsr/_0171_ ;
wire \mcsr/_0172_ ;
wire \mcsr/_0173_ ;
wire \mcsr/_0174_ ;
wire \mcsr/_0175_ ;
wire \mcsr/_0176_ ;
wire \mcsr/_0177_ ;
wire \mcsr/_0178_ ;
wire \mcsr/_0179_ ;
wire \mcsr/_0180_ ;
wire \mcsr/_0181_ ;
wire \mcsr/_0182_ ;
wire \mcsr/_0183_ ;
wire \mcsr/_0184_ ;
wire \mcsr/_0185_ ;
wire \mcsr/_0186_ ;
wire \mcsr/_0187_ ;
wire \mcsr/_0188_ ;
wire \mcsr/_0189_ ;
wire \mcsr/_0190_ ;
wire \mcsr/_0191_ ;
wire \mcsr/_0192_ ;
wire \mcsr/_0193_ ;
wire \mcsr/_0194_ ;
wire \mcsr/_0195_ ;
wire \mcsr/_0196_ ;
wire \mcsr/_0197_ ;
wire \mcsr/_0198_ ;
wire \mcsr/_0199_ ;
wire \mcsr/_0200_ ;
wire \mcsr/_0201_ ;
wire \mcsr/_0202_ ;
wire \mcsr/_0203_ ;
wire \mcsr/_0204_ ;
wire \mcsr/_0205_ ;
wire \mcsr/_0206_ ;
wire \mcsr/_0207_ ;
wire \mcsr/_0208_ ;
wire \mcsr/_0209_ ;
wire \mcsr/_0210_ ;
wire \mcsr/_0211_ ;
wire \mcsr/_0212_ ;
wire \mcsr/_0213_ ;
wire \mcsr/_0214_ ;
wire \mcsr/_0215_ ;
wire \mcsr/_0216_ ;
wire \mcsr/_0217_ ;
wire \mcsr/_0218_ ;
wire \mcsr/_0219_ ;
wire \mcsr/_0220_ ;
wire \mcsr/_0221_ ;
wire \mcsr/_0222_ ;
wire \mcsr/_0223_ ;
wire \mcsr/_0224_ ;
wire \mcsr/_0225_ ;
wire \mcsr/_0226_ ;
wire \mcsr/_0227_ ;
wire \mcsr/_0228_ ;
wire \mcsr/_0229_ ;
wire \mcsr/_0230_ ;
wire \mcsr/_0231_ ;
wire \mcsr/_0232_ ;
wire \mcsr/_0233_ ;
wire \mcsr/_0234_ ;
wire \mcsr/_0235_ ;
wire \mcsr/_0236_ ;
wire \mcsr/_0237_ ;
wire \mcsr/_0238_ ;
wire \mcsr/_0239_ ;
wire \mcsr/_0240_ ;
wire \mcsr/_0241_ ;
wire \mcsr/_0242_ ;
wire \mcsr/_0243_ ;
wire \mcsr/_0244_ ;
wire \mcsr/_0245_ ;
wire \mcsr/_0246_ ;
wire \mcsr/_0247_ ;
wire \mcsr/_0248_ ;
wire \mcsr/_0249_ ;
wire \mcsr/_0250_ ;
wire \mcsr/_0251_ ;
wire \mcsr/_0252_ ;
wire \mcsr/_0253_ ;
wire \mcsr/_0254_ ;
wire \mcsr/_0255_ ;
wire \mcsr/_0256_ ;
wire \mcsr/_0257_ ;
wire \mcsr/_0258_ ;
wire \mcsr/_0259_ ;
wire \mcsr/_0260_ ;
wire \mcsr/_0261_ ;
wire \mcsr/_0262_ ;
wire \mcsr/_0263_ ;
wire \mcsr/_0264_ ;
wire \mcsr/_0265_ ;
wire \mcsr/_0266_ ;
wire \mcsr/_0267_ ;
wire \mcsr/_0268_ ;
wire \mcsr/_0269_ ;
wire \mcsr/_0270_ ;
wire \mcsr/_0271_ ;
wire \mcsr/_0272_ ;
wire \mcsr/_0273_ ;
wire \mcsr/_0274_ ;
wire \mcsr/_0275_ ;
wire \mcsr/_0276_ ;
wire \mcsr/_0277_ ;
wire \mcsr/_0278_ ;
wire \mcsr/_0279_ ;
wire \mcsr/_0280_ ;
wire \mcsr/_0281_ ;
wire \mcsr/_0282_ ;
wire \mcsr/_0283_ ;
wire \mcsr/_0284_ ;
wire \mcsr/_0285_ ;
wire \mcsr/_0286_ ;
wire \mcsr/_0287_ ;
wire \mcsr/_0288_ ;
wire \mcsr/_0289_ ;
wire \mcsr/_0290_ ;
wire \mcsr/_0291_ ;
wire \mcsr/_0292_ ;
wire \mcsr/_0293_ ;
wire \mcsr/_0294_ ;
wire \mcsr/_0295_ ;
wire \mcsr/_0296_ ;
wire \mcsr/_0297_ ;
wire \mcsr/_0298_ ;
wire \mcsr/_0299_ ;
wire \mcsr/_0300_ ;
wire \mcsr/_0301_ ;
wire \mcsr/_0302_ ;
wire \mcsr/_0303_ ;
wire \mcsr/_0304_ ;
wire \mcsr/_0305_ ;
wire \mcsr/_0306_ ;
wire \mcsr/_0307_ ;
wire \mcsr/_0308_ ;
wire \mcsr/_0309_ ;
wire \mcsr/_0310_ ;
wire \mcsr/_0311_ ;
wire \mcsr/_0312_ ;
wire \mcsr/_0313_ ;
wire \mcsr/_0314_ ;
wire \mcsr/_0315_ ;
wire \mcsr/_0316_ ;
wire \mcsr/_0317_ ;
wire \mcsr/_0318_ ;
wire \mcsr/_0319_ ;
wire \mcsr/_0320_ ;
wire \mcsr/_0321_ ;
wire \mcsr/_0322_ ;
wire \mcsr/_0323_ ;
wire \mcsr/_0324_ ;
wire \mcsr/_0325_ ;
wire \mcsr/_0326_ ;
wire \mcsr/_0327_ ;
wire \mcsr/_0328_ ;
wire \mcsr/_0329_ ;
wire \mcsr/_0330_ ;
wire \mcsr/_0331_ ;
wire \mcsr/_0332_ ;
wire \mcsr/_0333_ ;
wire \mcsr/_0334_ ;
wire \mcsr/_0335_ ;
wire \mcsr/_0336_ ;
wire \mcsr/_0337_ ;
wire \mcsr/_0338_ ;
wire \mcsr/_0339_ ;
wire \mcsr/_0340_ ;
wire \mcsr/_0341_ ;
wire \mcsr/_0342_ ;
wire \mcsr/_0343_ ;
wire \mcsr/_0344_ ;
wire \mcsr/_0345_ ;
wire \mcsr/_0346_ ;
wire \mcsr/_0347_ ;
wire \mcsr/_0348_ ;
wire \mcsr/_0349_ ;
wire \mcsr/_0350_ ;
wire \mcsr/_0351_ ;
wire \mcsr/_0352_ ;
wire \mcsr/_0353_ ;
wire \mcsr/_0354_ ;
wire \mcsr/_0355_ ;
wire \mcsr/_0356_ ;
wire \mcsr/_0357_ ;
wire \mcsr/_0358_ ;
wire \mcsr/_0359_ ;
wire \mcsr/_0360_ ;
wire \mcsr/_0361_ ;
wire \mcsr/_0362_ ;
wire \mcsr/_0363_ ;
wire \mcsr/_0364_ ;
wire \mcsr/_0365_ ;
wire \mcsr/_0366_ ;
wire \mcsr/_0367_ ;
wire \mcsr/_0368_ ;
wire \mcsr/_0369_ ;
wire \mcsr/_0370_ ;
wire \mcsr/_0371_ ;
wire \mcsr/_0372_ ;
wire \mcsr/_0373_ ;
wire \mcsr/_0374_ ;
wire \mcsr/_0375_ ;
wire \mcsr/_0376_ ;
wire \mcsr/_0377_ ;
wire \mcsr/_0378_ ;
wire \mcsr/_0379_ ;
wire \mcsr/_0380_ ;
wire \mcsr/_0381_ ;
wire \mcsr/_0382_ ;
wire \mcsr/_0383_ ;
wire \mcsr/_0384_ ;
wire \mcsr/_0385_ ;
wire \mcsr/_0386_ ;
wire \mcsr/_0387_ ;
wire \mcsr/_0388_ ;
wire \mcsr/_0389_ ;
wire \mcsr/_0390_ ;
wire \mcsr/_0391_ ;
wire \mcsr/_0392_ ;
wire \mcsr/_0393_ ;
wire \mcsr/_0394_ ;
wire \mcsr/_0395_ ;
wire \mcsr/_0396_ ;
wire \mcsr/_0397_ ;
wire \mcsr/_0398_ ;
wire \mcsr/_0399_ ;
wire \mcsr/_0400_ ;
wire \mcsr/_0401_ ;
wire \mcsr/_0402_ ;
wire \mcsr/_0403_ ;
wire \mcsr/_0404_ ;
wire \mcsr/_0405_ ;
wire \mcsr/_0406_ ;
wire \mcsr/_0407_ ;
wire \mcsr/_0408_ ;
wire \mcsr/_0409_ ;
wire \mcsr/_0410_ ;
wire \mcsr/_0411_ ;
wire \mcsr/_0412_ ;
wire \mcsr/_0413_ ;
wire \mcsr/_0414_ ;
wire \mcsr/_0415_ ;
wire \mcsr/_0416_ ;
wire \mcsr/_0417_ ;
wire \mcsr/_0418_ ;
wire \mcsr/_0419_ ;
wire \mcsr/_0420_ ;
wire \mcsr/_0421_ ;
wire \mcsr/_0422_ ;
wire \mcsr/_0423_ ;
wire \mcsr/_0424_ ;
wire \mcsr/_0425_ ;
wire \mcsr/_0426_ ;
wire \mcsr/_0427_ ;
wire \mcsr/_0428_ ;
wire \mcsr/_0429_ ;
wire \mcsr/_0430_ ;
wire \mcsr/_0431_ ;
wire \mcsr/_0432_ ;
wire \mcsr/_0433_ ;
wire \mcsr/_0434_ ;
wire \mcsr/_0435_ ;
wire \mcsr/_0436_ ;
wire \mcsr/_0437_ ;
wire \mcsr/_0438_ ;
wire \mcsr/_0439_ ;
wire \mcsr/_0440_ ;
wire \mcsr/_0441_ ;
wire \mcsr/_0442_ ;
wire \mcsr/_0443_ ;
wire \mcsr/_0444_ ;
wire \mcsr/_0445_ ;
wire \mcsr/_0446_ ;
wire \mcsr/_0447_ ;
wire \mcsr/_0448_ ;
wire \mcsr/_0449_ ;
wire \mcsr/_0450_ ;
wire \mcsr/_0451_ ;
wire \mcsr/_0452_ ;
wire \mcsr/_0453_ ;
wire \mcsr/_0454_ ;
wire \mcsr/_0455_ ;
wire \mcsr/_0456_ ;
wire \mcsr/_0457_ ;
wire \mcsr/_0458_ ;
wire \mcsr/_0459_ ;
wire \mcsr/_0460_ ;
wire \mcsr/_0461_ ;
wire \mcsr/_0462_ ;
wire \mcsr/_0463_ ;
wire \mcsr/_0464_ ;
wire \mcsr/_0465_ ;
wire \mcsr/_0466_ ;
wire \mcsr/_0467_ ;
wire \mcsr/_0468_ ;
wire \mcsr/_0469_ ;
wire \mcsr/_0470_ ;
wire \mcsr/_0471_ ;
wire \mcsr/_0472_ ;
wire \mcsr/_0473_ ;
wire \mcsr/_0474_ ;
wire \mcsr/_0475_ ;
wire \mcsr/_0476_ ;
wire \mcsr/_0477_ ;
wire \mcsr/_0478_ ;
wire \mcsr/_0479_ ;
wire \mcsr/_0480_ ;
wire \mcsr/_0481_ ;
wire \mcsr/_0482_ ;
wire \mcsr/_0483_ ;
wire \mcsr/_0484_ ;
wire \mcsr/_0485_ ;
wire \mcsr/_0486_ ;
wire \mcsr/_0487_ ;
wire \mcsr/_0488_ ;
wire \mcsr/_0489_ ;
wire \mcsr/_0490_ ;
wire \mcsr/_0491_ ;
wire \mcsr/_0492_ ;
wire \mcsr/_0493_ ;
wire \mcsr/_0494_ ;
wire \mcsr/_0495_ ;
wire \mcsr/_0496_ ;
wire \mcsr/_0497_ ;
wire \mcsr/_0498_ ;
wire \mcsr/_0499_ ;
wire \mcsr/_0500_ ;
wire \mcsr/_0501_ ;
wire \mcsr/_0502_ ;
wire \mcsr/_0503_ ;
wire \mcsr/_0504_ ;
wire \mcsr/_0505_ ;
wire \mcsr/_0506_ ;
wire \mcsr/_0507_ ;
wire \mcsr/_0508_ ;
wire \mcsr/_0509_ ;
wire \mcsr/_0510_ ;
wire \mcsr/_0511_ ;
wire \mcsr/_0512_ ;
wire \mcsr/_0513_ ;
wire \mcsr/_0514_ ;
wire \mcsr/_0515_ ;
wire \mcsr/_0516_ ;
wire \mcsr/_0517_ ;
wire \mcsr/_0518_ ;
wire \mcsr/_0519_ ;
wire \mcsr/_0520_ ;
wire \mcsr/_0521_ ;
wire \mcsr/_0522_ ;
wire \mcsr/_0523_ ;
wire \mcsr/_0524_ ;
wire \mcsr/_0525_ ;
wire \mcsr/_0526_ ;
wire \mcsr/_0527_ ;
wire \mcsr/_0528_ ;
wire \mcsr/_0529_ ;
wire \mcsr/_0530_ ;
wire \mcsr/_0531_ ;
wire \mcsr/_0532_ ;
wire \mcsr/_0533_ ;
wire \mcsr/_0534_ ;
wire \mcsr/_0535_ ;
wire \mcsr/_0536_ ;
wire \mcsr/_0537_ ;
wire \mcsr/_0538_ ;
wire \mcsr/_0539_ ;
wire \mcsr/_0540_ ;
wire \mcsr/_0541_ ;
wire \mcsr/_0542_ ;
wire \mcsr/_0543_ ;
wire \mcsr/_0544_ ;
wire \mcsr/_0545_ ;
wire \mcsr/_0546_ ;
wire \mcsr/_0547_ ;
wire \mcsr/_0548_ ;
wire \mcsr/_0549_ ;
wire \mcsr/_0550_ ;
wire \mcsr/_0551_ ;
wire \mcsr/_0552_ ;
wire \mcsr/_0553_ ;
wire \mcsr/_0554_ ;
wire \mcsr/_0555_ ;
wire \mcsr/_0556_ ;
wire \mcsr/_0557_ ;
wire \mcsr/_0558_ ;
wire \mcsr/_0559_ ;
wire \mcsr/_0560_ ;
wire \mcsr/_0561_ ;
wire \mcsr/_0562_ ;
wire \mcsr/_0563_ ;
wire \mcsr/_0564_ ;
wire \mcsr/_0565_ ;
wire \mcsr/_0566_ ;
wire \mcsr/_0567_ ;
wire \mcsr/_0568_ ;
wire \mcsr/_0569_ ;
wire \mcsr/_0570_ ;
wire \mcsr/_0571_ ;
wire \mcsr/_0572_ ;
wire \mcsr/_0573_ ;
wire \mcsr/_0574_ ;
wire \mcsr/_0575_ ;
wire \mcsr/_0576_ ;
wire \mcsr/_0577_ ;
wire \mcsr/_0578_ ;
wire \mcsr/_0579_ ;
wire \mcsr/_0580_ ;
wire \mcsr/_0581_ ;
wire \mcsr/_0582_ ;
wire \mcsr/_0583_ ;
wire \mcsr/_0584_ ;
wire \mcsr/_0585_ ;
wire \mcsr/_0586_ ;
wire \mcsr/_0587_ ;
wire \mcsr/_0588_ ;
wire \mcsr/_0589_ ;
wire \mcsr/_0590_ ;
wire \mcsr/_0591_ ;
wire \mcsr/_0592_ ;
wire \mcsr/_0593_ ;
wire \mcsr/_0594_ ;
wire \mcsr/_0595_ ;
wire \mcsr/_0596_ ;
wire \mcsr/_0597_ ;
wire \mcsr/_0598_ ;
wire \mcsr/_0599_ ;
wire \mcsr/_0600_ ;
wire \mcsr/_0601_ ;
wire \mcsr/_0602_ ;
wire \mcsr/_0603_ ;
wire \mcsr/_0604_ ;
wire \mcsr/_0605_ ;
wire \mcsr/_0606_ ;
wire \mcsr/_0607_ ;
wire \mcsr/_0608_ ;
wire \mcsr/_0609_ ;
wire \mcsr/_0610_ ;
wire \mcsr/_0611_ ;
wire \mcsr/_0612_ ;
wire \mcsr/_0613_ ;
wire \mcsr/_0614_ ;
wire \mcsr/_0615_ ;
wire \mcsr/_0616_ ;
wire \mcsr/_0617_ ;
wire \mcsr/_0618_ ;
wire \mcsr/_0619_ ;
wire \mcsr/_0620_ ;
wire \mcsr/_0621_ ;
wire \mcsr/_0622_ ;
wire \mcsr/_0623_ ;
wire \mcsr/_0624_ ;
wire \mcsr/_0625_ ;
wire \mcsr/_0626_ ;
wire \mcsr/_0627_ ;
wire \mcsr/_0628_ ;
wire \mcsr/_0629_ ;
wire \mcsr/_0630_ ;
wire \mcsr/_0631_ ;
wire \mcsr/_0632_ ;
wire \mcsr/_0633_ ;
wire \mcsr/_0634_ ;
wire \mcsr/_0635_ ;
wire \mcsr/_0636_ ;
wire \mcsr/_0637_ ;
wire \mcsr/_0638_ ;
wire \mcsr/_0639_ ;
wire \mcsr/_0640_ ;
wire \mcsr/_0641_ ;
wire \mcsr/_0642_ ;
wire \mcsr/_0643_ ;
wire \mcsr/_0644_ ;
wire \mcsr/_0645_ ;
wire \mcsr/_0646_ ;
wire \mcsr/_0647_ ;
wire \mcsr/_0648_ ;
wire \mcsr/_0649_ ;
wire \mcsr/_0650_ ;
wire \mcsr/_0651_ ;
wire \mcsr/_0652_ ;
wire \mcsr/_0653_ ;
wire \mcsr/_0654_ ;
wire \mcsr/_0655_ ;
wire \mcsr/_0656_ ;
wire \mcsr/_0657_ ;
wire \mcsr/_0658_ ;
wire \mcsr/_0659_ ;
wire \mcsr/_0660_ ;
wire \mcsr/_0661_ ;
wire \mcsr/_0662_ ;
wire \mcsr/_0663_ ;
wire \mcsr/_0664_ ;
wire \mcsr/_0665_ ;
wire \mcsr/_0666_ ;
wire \mcsr/_0667_ ;
wire \mcsr/_0668_ ;
wire \mcsr/_0669_ ;
wire \mcsr/_0670_ ;
wire \mcsr/_0671_ ;
wire \mcsr/_0672_ ;
wire \mcsr/_0673_ ;
wire \mcsr/_0674_ ;
wire \mcsr/_0675_ ;
wire \mcsr/_0676_ ;
wire \mcsr/_0677_ ;
wire \mcsr/_0678_ ;
wire \mcsr/_0679_ ;
wire \mcsr/_0680_ ;
wire \mcsr/_0681_ ;
wire \mcsr/_0682_ ;
wire \mcsr/_0683_ ;
wire \mcsr/_0684_ ;
wire \mcsr/_0685_ ;
wire \mcsr/_0686_ ;
wire \mcsr/_0687_ ;
wire \mcsr/_0688_ ;
wire \mcsr/_0689_ ;
wire \mcsr/_0690_ ;
wire \mcsr/_0691_ ;
wire \mcsr/_0692_ ;
wire \mcsr/_0693_ ;
wire \mcsr/_0694_ ;
wire \mcsr/_0695_ ;
wire \mcsr/_0696_ ;
wire \mcsr/_0697_ ;
wire \mcsr/_0698_ ;
wire \mcsr/_0699_ ;
wire \mcsr/_0700_ ;
wire \mcsr/_0701_ ;
wire \mcsr/_0702_ ;
wire \mcsr/_0703_ ;
wire \mcsr/_0704_ ;
wire \mcsr/_0705_ ;
wire \mcsr/_0706_ ;
wire \mcsr/_0707_ ;
wire \mcsr/_0708_ ;
wire \mcsr/_0709_ ;
wire \mcsr/_0710_ ;
wire \mcsr/_0711_ ;
wire \mcsr/_0712_ ;
wire \mcsr/_0713_ ;
wire \mcsr/_0714_ ;
wire \mcsr/_0715_ ;
wire \mcsr/_0716_ ;
wire \mcsr/_0717_ ;
wire \mcsr/_0718_ ;
wire \mcsr/_0719_ ;
wire \mcsr/_0720_ ;
wire \mcsr/_0721_ ;
wire \mcsr/_0722_ ;
wire \mcsr/_0723_ ;
wire \mcsr/_0724_ ;
wire \mcsr/_0725_ ;
wire \mcsr/_0726_ ;
wire \mcsr/_0727_ ;
wire \mcsr/_0728_ ;
wire \mcsr/_0729_ ;
wire \mcsr/_0730_ ;
wire \mcsr/_0731_ ;
wire \mcsr/_0732_ ;
wire \mcsr/_0733_ ;
wire \mcsr/_0734_ ;
wire \mcsr/_0735_ ;
wire \mcsr/_0736_ ;
wire \mcsr/_0737_ ;
wire \mcsr/_0738_ ;
wire \mcsr/_0739_ ;
wire \mcsr/_0740_ ;
wire \mcsr/_0741_ ;
wire \mcsr/_0742_ ;
wire \mcsr/_0743_ ;
wire \mcsr/_0744_ ;
wire \mcsr/_0745_ ;
wire \mcsr/_0746_ ;
wire \mcsr/_0747_ ;
wire \mcsr/_0748_ ;
wire \mcsr/_0749_ ;
wire \mcsr/_0750_ ;
wire \mcsr/_0751_ ;
wire \mcsr/_0752_ ;
wire \mcsr/_0753_ ;
wire \mcsr/_0754_ ;
wire \mcsr/_0755_ ;
wire \mcsr/_0756_ ;
wire \mcsr/_0757_ ;
wire \mcsr/_0758_ ;
wire \mcsr/_0759_ ;
wire \mcsr/_0760_ ;
wire \mcsr/_0761_ ;
wire \mcsr/_0762_ ;
wire \mcsr/_0763_ ;
wire \mcsr/_0764_ ;
wire \mcsr/_0765_ ;
wire \mcsr/_0766_ ;
wire \mcsr/_0767_ ;
wire \mcsr/_0768_ ;
wire \mcsr/_0769_ ;
wire \mcsr/_0770_ ;
wire \mcsr/_0771_ ;
wire \mcsr/_0772_ ;
wire \mcsr/_0773_ ;
wire \mcsr/_0774_ ;
wire \mcsr/_0775_ ;
wire \mcsr/_0776_ ;
wire \mcsr/_0777_ ;
wire \mcsr/_0778_ ;
wire \mcsr/_0779_ ;
wire \mcsr/_0780_ ;
wire \mcsr/_0781_ ;
wire \mcsr/_0782_ ;
wire \mcsr/_0783_ ;
wire \mcsr/_0784_ ;
wire \mcsr/_0785_ ;
wire \mcsr/_0786_ ;
wire \mcsr/_0787_ ;
wire \mcsr/_0788_ ;
wire \mcsr/_0789_ ;
wire \mcsr/_0790_ ;
wire \mcsr/_0791_ ;
wire \mcsr/_0792_ ;
wire \mcsr/_0793_ ;
wire \mcsr/_0794_ ;
wire \mcsr/_0795_ ;
wire \mcsr/_0796_ ;
wire \mcsr/_0797_ ;
wire \mcsr/_0798_ ;
wire \mcsr/_0799_ ;
wire \mcsr/_0800_ ;
wire \mcsr/_0801_ ;
wire \mcsr/_0802_ ;
wire \mcsr/_0803_ ;
wire \mcsr/_0804_ ;
wire \mcsr/_0805_ ;
wire \mcsr/_0806_ ;
wire \mcsr/_0807_ ;
wire \mcsr/_0808_ ;
wire \mcsr/_0809_ ;
wire \mcsr/_0810_ ;
wire \mcsr/_0811_ ;
wire \mcsr/_0812_ ;
wire \mcsr/_0813_ ;
wire \mcsr/_0814_ ;
wire \mcsr/_0815_ ;
wire \mcsr/_0816_ ;
wire \mcsr/_0817_ ;
wire \mcsr/_0818_ ;
wire \mcsr/_0819_ ;
wire \mcsr/_0820_ ;
wire \mcsr/_0821_ ;
wire \mcsr/_0822_ ;
wire \mcsr/_0823_ ;
wire \mcsr/_0824_ ;
wire \mcsr/_0825_ ;
wire \mcsr/_0826_ ;
wire \mcsr/_0827_ ;
wire \mcsr/_0828_ ;
wire \mcsr/_0829_ ;
wire \mcsr/_0830_ ;
wire \mcsr/_0831_ ;
wire \mcsr/_0832_ ;
wire \mcsr/_0833_ ;
wire \mcsr/_0834_ ;
wire \mcsr/_0835_ ;
wire \mcsr/_0836_ ;
wire \mcsr/_0837_ ;
wire \mcsr/_0838_ ;
wire \mcsr/_0839_ ;
wire \mcsr/_0840_ ;
wire \mcsr/_0841_ ;
wire \mcsr/_0842_ ;
wire \mcsr/_0843_ ;
wire \mcsr/_0844_ ;
wire \mcsr/_0845_ ;
wire \mcsr/_0846_ ;
wire \mcsr/_0847_ ;
wire \mcsr/_0848_ ;
wire \mcsr/_0849_ ;
wire \mcsr/_0850_ ;
wire \mcsr/_0851_ ;
wire \mcsr/_0852_ ;
wire \mcsr/_0853_ ;
wire \mcsr/_0854_ ;
wire \mcsr/_0855_ ;
wire \mcsr/_0856_ ;
wire \mcsr/_0857_ ;
wire \mcsr/_0858_ ;
wire \mcsr/_0859_ ;
wire \mcsr/_0860_ ;
wire \mcsr/_0861_ ;
wire \mcsr/_0862_ ;
wire \mcsr/_0863_ ;
wire \mcsr/_0864_ ;
wire \mcsr/_0865_ ;
wire \mcsr/_0866_ ;
wire \mcsr/_0867_ ;
wire \mcsr/_0868_ ;
wire \mcsr/_0869_ ;
wire \mcsr/_0870_ ;
wire \mcsr/_0871_ ;
wire \mcsr/_0872_ ;
wire \mcsr/_0873_ ;
wire \mcsr/_0874_ ;
wire \mcsr/_0875_ ;
wire \mcsr/_0876_ ;
wire \mcsr/_0877_ ;
wire \mcsr/_0878_ ;
wire \mcsr/_0879_ ;
wire \mcsr/_0880_ ;
wire \mcsr/_0881_ ;
wire \mcsr/_0882_ ;
wire \mcsr/_0883_ ;
wire \mcsr/_0884_ ;
wire \mcsr/_0885_ ;
wire \mcsr/_0886_ ;
wire \mcsr/_0887_ ;
wire \mcsr/_0888_ ;
wire \mcsr/_0889_ ;
wire \mcsr/_0890_ ;
wire \mcsr/_0891_ ;
wire \mcsr/_0892_ ;
wire \mcsr/_0893_ ;
wire \mcsr/_0894_ ;
wire \mcsr/_0895_ ;
wire \mcsr/_0896_ ;
wire \mcsr/_0897_ ;
wire \mcsr/_0898_ ;
wire \mcsr/_0899_ ;
wire \mcsr/_0900_ ;
wire \mcsr/_0901_ ;
wire \mcsr/_0902_ ;
wire \mcsr/_0903_ ;
wire \mcsr/_0904_ ;
wire \mcsr/_0905_ ;
wire \mcsr/_0906_ ;
wire \mcsr/_0907_ ;
wire \mcsr/_0908_ ;
wire \mcsr/_0909_ ;
wire \mcsr/_0910_ ;
wire \mcsr/_0911_ ;
wire \mcsr/_0912_ ;
wire \mcsr/_0913_ ;
wire \mcsr/_0914_ ;
wire \mcsr/_0915_ ;
wire \mcsr/_0916_ ;
wire \mcsr/_0917_ ;
wire \mcsr/_0918_ ;
wire \mcsr/_0919_ ;
wire \mcsr/_0920_ ;
wire \mcsr/_0921_ ;
wire \mcsr/_0922_ ;
wire \mcsr/_0923_ ;
wire \mcsr/_0924_ ;
wire \mcsr/_0925_ ;
wire \mcsr/_0926_ ;
wire \mcsr/_0927_ ;
wire \mcsr/_0928_ ;
wire \mcsr/_0929_ ;
wire \mcsr/_0930_ ;
wire \mcsr/_0931_ ;
wire \mcsr/_0932_ ;
wire \mcsr/_0933_ ;
wire \mcsr/_0934_ ;
wire \mcsr/_0935_ ;
wire \mcsr/_0936_ ;
wire \mcsr/_0937_ ;
wire \mcsr/_0938_ ;
wire \mcsr/_0939_ ;
wire \mcsr/_0940_ ;
wire \mcsr/_0941_ ;
wire \mcsr/_0942_ ;
wire \mcsr/_0943_ ;
wire \mcsr/_0944_ ;
wire \mcsr/_0945_ ;
wire \mcsr/_0946_ ;
wire \mcsr/_0947_ ;
wire \mcsr/_0948_ ;
wire \mcsr/_0949_ ;
wire \mcsr/_0950_ ;
wire \mcsr/_0951_ ;
wire \mcsr/_0952_ ;
wire \mcsr/_0953_ ;
wire \mcsr/_0954_ ;
wire \mcsr/_0955_ ;
wire \mcsr/_0956_ ;
wire \mcsr/_0957_ ;
wire \mcsr/_0958_ ;
wire \mcsr/_0959_ ;
wire \mcsr/_0960_ ;
wire \mcsr/_0961_ ;
wire \mcsr/_0962_ ;
wire \mcsr/_0963_ ;
wire \mcsr/_0964_ ;
wire \mcsr/_0965_ ;
wire \mcsr/_0966_ ;
wire \mcsr/_0967_ ;
wire \mcsr/_0968_ ;
wire \mcsr/_0969_ ;
wire \mcsr/_0970_ ;
wire \mcsr/_0971_ ;
wire \mcsr/_0972_ ;
wire \mcsr/_0973_ ;
wire \mcsr/_0974_ ;
wire \mcsr/_0975_ ;
wire \mcsr/_0976_ ;
wire \mcsr/_0977_ ;
wire \mcsr/_0978_ ;
wire \mcsr/_0979_ ;
wire \mcsr/_0980_ ;
wire \mcsr/_0981_ ;
wire \mcsr/_0982_ ;
wire \mcsr/_0983_ ;
wire \mcsr/_0984_ ;
wire \mcsr/_0985_ ;
wire \mcsr/_0986_ ;
wire \mcsr/_0987_ ;
wire \mcsr/_0988_ ;
wire \mcsr/_0989_ ;
wire \mcsr/_0990_ ;
wire \mcsr/_0991_ ;
wire \mcsr/_0992_ ;
wire \mcsr/_0993_ ;
wire \mcsr/_0994_ ;
wire \mcsr/_0995_ ;
wire \mcsr/_0996_ ;
wire \mcsr/_0997_ ;
wire \mcsr/_0998_ ;
wire \mcsr/_0999_ ;
wire \mcsr/_1000_ ;
wire \mcsr/_1001_ ;
wire \mcsr/_1002_ ;
wire \mcsr/_1003_ ;
wire \mcsr/_1004_ ;
wire \mcsr/_1005_ ;
wire \mcsr/_1006_ ;
wire \mcsr/_1007_ ;
wire \mcsr/_1008_ ;
wire \mcsr/_1009_ ;
wire \mcsr/_1010_ ;
wire \mcsr/_1011_ ;
wire \mcsr/_1012_ ;
wire \mcsr/_1013_ ;
wire \mcsr/_1014_ ;
wire \mcsr/_1015_ ;
wire \mcsr/_1016_ ;
wire \mcsr/_1017_ ;
wire \mcsr/_1018_ ;
wire \mcsr/_1019_ ;
wire \mcsr/_1020_ ;
wire \mcsr/_1021_ ;
wire \mcsr/_1022_ ;
wire \mcsr/_1023_ ;
wire \mcsr/_1024_ ;
wire \mcsr/_1025_ ;
wire \mcsr/_1026_ ;
wire \mcsr/_1027_ ;
wire \mcsr/_1028_ ;
wire \mcsr/_1029_ ;
wire \mcsr/_1030_ ;
wire \mcsr/_1031_ ;
wire \mcsr/_1032_ ;
wire \mcsr/_1033_ ;
wire \mcsr/_1034_ ;
wire \mcsr/_1035_ ;
wire \mcsr/_1036_ ;
wire \mcsr/_1037_ ;
wire \mcsr/_1038_ ;
wire \mcsr/_1039_ ;
wire \mcsr/_1040_ ;
wire \mcsr/_1041_ ;
wire \mcsr/_1042_ ;
wire \mcsr/_1043_ ;
wire \mcsr/_1044_ ;
wire \mcsr/_1045_ ;
wire \mcsr/_1046_ ;
wire \mcsr/_1047_ ;
wire \mcsr/_1048_ ;
wire \mcsr/_1049_ ;
wire \mcsr/_1050_ ;
wire \mcsr/_1051_ ;
wire \mcsr/_1052_ ;
wire \mcsr/_1053_ ;
wire \mcsr/_1054_ ;
wire \mcsr/_1055_ ;
wire \mcsr/_1056_ ;
wire \mcsr/_1057_ ;
wire \mcsr/_1058_ ;
wire \mcsr/_1059_ ;
wire \mcsr/_1060_ ;
wire \mcsr/_1061_ ;
wire \mcsr/_1062_ ;
wire \mcsr/_1063_ ;
wire \mcsr/_1064_ ;
wire \mcsr/_1065_ ;
wire \mcsr/_1066_ ;
wire \mcsr/_1067_ ;
wire \mcsr/_1068_ ;
wire \mcsr/_1069_ ;
wire \mcsr/_1070_ ;
wire \mcsr/_1071_ ;
wire \mcsr/_1072_ ;
wire \mcsr/_1073_ ;
wire \mcsr/_1074_ ;
wire \mcsr/_1075_ ;
wire \mcsr/_1076_ ;
wire \mcsr/_1077_ ;
wire \mcsr/_1078_ ;
wire \mcsr/_1079_ ;
wire \mcsr/_1080_ ;
wire \mcsr/_1081_ ;
wire \mcsr/_1082_ ;
wire \mcsr/_1083_ ;
wire \mcsr/_1084_ ;
wire \mcsr/_1085_ ;
wire \mcsr/_1086_ ;
wire \mcsr/_1087_ ;
wire \mcsr/_1088_ ;
wire \mcsr/_1089_ ;
wire \mcsr/_1090_ ;
wire \mcsr/_1091_ ;
wire \mcsr/_1092_ ;
wire \mcsr/_1093_ ;
wire \mcsr/_1094_ ;
wire \mcsr/_1095_ ;
wire \mcsr/_1096_ ;
wire \mcsr/_1097_ ;
wire \mcsr/_1098_ ;
wire \mcsr/_1099_ ;
wire \mcsr/_1100_ ;
wire \mcsr/_1101_ ;
wire \mcsr/_1102_ ;
wire \mcsr/_1103_ ;
wire \mcsr/_1104_ ;
wire \mcsr/_1105_ ;
wire \mcsr/_1106_ ;
wire \mcsr/_1107_ ;
wire \mcsr/_1108_ ;
wire \mcsr/_1109_ ;
wire \mcsr/_1110_ ;
wire \mcsr/_1111_ ;
wire \mcsr/_1112_ ;
wire \mcsr/_1113_ ;
wire \mcsr/_1114_ ;
wire \mcsr/_1115_ ;
wire \mcsr/_1116_ ;
wire \mcsr/_1117_ ;
wire \mcsr/_1118_ ;
wire \mcsr/_1119_ ;
wire \mcsr/_1120_ ;
wire \mcsr/_1121_ ;
wire \mcsr/_1122_ ;
wire \mcsr/_1123_ ;
wire \mcsr/_1124_ ;
wire \mcsr/_1125_ ;
wire \mcsr/_1126_ ;
wire \mcsr/_1127_ ;
wire \mcsr/_1128_ ;
wire \mcsr/_1129_ ;
wire \mcsr/_1130_ ;
wire \mcsr/_1131_ ;
wire \mcsr/_1132_ ;
wire \mcsr/_1133_ ;
wire \mcsr/_1134_ ;
wire \mcsr/_1135_ ;
wire \mcsr/_1136_ ;
wire \mcsr/_1137_ ;
wire \mcsr/_1138_ ;
wire \mcsr/_1139_ ;
wire \mcsr/_1140_ ;
wire \mcsr/_1141_ ;
wire \mcsr/_1142_ ;
wire \mcsr/_1143_ ;
wire \mcsr/_1144_ ;
wire \mcsr/_1145_ ;
wire \mcsr/_1146_ ;
wire \mcsr/_1147_ ;
wire \mcsr/_1148_ ;
wire \mcsr/_1149_ ;
wire \mcsr/_1150_ ;
wire \mcsr/_1151_ ;
wire \mcsr/_1152_ ;
wire \mcsr/_1153_ ;
wire \mcsr/_1154_ ;
wire \mcsr/csr[0][0] ;
wire \mcsr/csr[0][10] ;
wire \mcsr/csr[0][11] ;
wire \mcsr/csr[0][12] ;
wire \mcsr/csr[0][13] ;
wire \mcsr/csr[0][14] ;
wire \mcsr/csr[0][15] ;
wire \mcsr/csr[0][16] ;
wire \mcsr/csr[0][17] ;
wire \mcsr/csr[0][18] ;
wire \mcsr/csr[0][19] ;
wire \mcsr/csr[0][1] ;
wire \mcsr/csr[0][20] ;
wire \mcsr/csr[0][21] ;
wire \mcsr/csr[0][22] ;
wire \mcsr/csr[0][23] ;
wire \mcsr/csr[0][24] ;
wire \mcsr/csr[0][25] ;
wire \mcsr/csr[0][26] ;
wire \mcsr/csr[0][27] ;
wire \mcsr/csr[0][28] ;
wire \mcsr/csr[0][29] ;
wire \mcsr/csr[0][2] ;
wire \mcsr/csr[0][30] ;
wire \mcsr/csr[0][31] ;
wire \mcsr/csr[0][3] ;
wire \mcsr/csr[0][4] ;
wire \mcsr/csr[0][5] ;
wire \mcsr/csr[0][6] ;
wire \mcsr/csr[0][7] ;
wire \mcsr/csr[0][8] ;
wire \mcsr/csr[0][9] ;
wire \mcsr/csr[1][0] ;
wire \mcsr/csr[1][10] ;
wire \mcsr/csr[1][11] ;
wire \mcsr/csr[1][12] ;
wire \mcsr/csr[1][13] ;
wire \mcsr/csr[1][14] ;
wire \mcsr/csr[1][15] ;
wire \mcsr/csr[1][16] ;
wire \mcsr/csr[1][17] ;
wire \mcsr/csr[1][18] ;
wire \mcsr/csr[1][19] ;
wire \mcsr/csr[1][1] ;
wire \mcsr/csr[1][20] ;
wire \mcsr/csr[1][21] ;
wire \mcsr/csr[1][22] ;
wire \mcsr/csr[1][23] ;
wire \mcsr/csr[1][24] ;
wire \mcsr/csr[1][25] ;
wire \mcsr/csr[1][26] ;
wire \mcsr/csr[1][27] ;
wire \mcsr/csr[1][28] ;
wire \mcsr/csr[1][29] ;
wire \mcsr/csr[1][2] ;
wire \mcsr/csr[1][30] ;
wire \mcsr/csr[1][31] ;
wire \mcsr/csr[1][3] ;
wire \mcsr/csr[1][4] ;
wire \mcsr/csr[1][5] ;
wire \mcsr/csr[1][6] ;
wire \mcsr/csr[1][7] ;
wire \mcsr/csr[1][8] ;
wire \mcsr/csr[1][9] ;
wire \mcsr/csr[2][0] ;
wire \mcsr/csr[2][10] ;
wire \mcsr/csr[2][11] ;
wire \mcsr/csr[2][12] ;
wire \mcsr/csr[2][13] ;
wire \mcsr/csr[2][14] ;
wire \mcsr/csr[2][15] ;
wire \mcsr/csr[2][16] ;
wire \mcsr/csr[2][17] ;
wire \mcsr/csr[2][18] ;
wire \mcsr/csr[2][19] ;
wire \mcsr/csr[2][1] ;
wire \mcsr/csr[2][20] ;
wire \mcsr/csr[2][21] ;
wire \mcsr/csr[2][22] ;
wire \mcsr/csr[2][23] ;
wire \mcsr/csr[2][24] ;
wire \mcsr/csr[2][25] ;
wire \mcsr/csr[2][26] ;
wire \mcsr/csr[2][27] ;
wire \mcsr/csr[2][28] ;
wire \mcsr/csr[2][29] ;
wire \mcsr/csr[2][2] ;
wire \mcsr/csr[2][30] ;
wire \mcsr/csr[2][31] ;
wire \mcsr/csr[2][3] ;
wire \mcsr/csr[2][4] ;
wire \mcsr/csr[2][5] ;
wire \mcsr/csr[2][6] ;
wire \mcsr/csr[2][7] ;
wire \mcsr/csr[2][8] ;
wire \mcsr/csr[2][9] ;
wire \mcsr/csr[3][0] ;
wire \mcsr/csr[3][10] ;
wire \mcsr/csr[3][11] ;
wire \mcsr/csr[3][12] ;
wire \mcsr/csr[3][13] ;
wire \mcsr/csr[3][14] ;
wire \mcsr/csr[3][15] ;
wire \mcsr/csr[3][16] ;
wire \mcsr/csr[3][17] ;
wire \mcsr/csr[3][18] ;
wire \mcsr/csr[3][19] ;
wire \mcsr/csr[3][1] ;
wire \mcsr/csr[3][20] ;
wire \mcsr/csr[3][21] ;
wire \mcsr/csr[3][22] ;
wire \mcsr/csr[3][23] ;
wire \mcsr/csr[3][24] ;
wire \mcsr/csr[3][25] ;
wire \mcsr/csr[3][26] ;
wire \mcsr/csr[3][27] ;
wire \mcsr/csr[3][28] ;
wire \mcsr/csr[3][29] ;
wire \mcsr/csr[3][2] ;
wire \mcsr/csr[3][30] ;
wire \mcsr/csr[3][31] ;
wire \mcsr/csr[3][3] ;
wire \mcsr/csr[3][4] ;
wire \mcsr/csr[3][5] ;
wire \mcsr/csr[3][6] ;
wire \mcsr/csr[3][7] ;
wire \mcsr/csr[3][8] ;
wire \mcsr/csr[3][9] ;
wire \mexu/_0000_ ;
wire \mexu/_0001_ ;
wire \mexu/_0002_ ;
wire \mexu/_0003_ ;
wire \mexu/_0004_ ;
wire \mexu/_0005_ ;
wire \mexu/_0006_ ;
wire \mexu/_0007_ ;
wire \mexu/_0008_ ;
wire \mexu/_0009_ ;
wire \mexu/_0010_ ;
wire \mexu/_0011_ ;
wire \mexu/_0012_ ;
wire \mexu/_0013_ ;
wire \mexu/_0014_ ;
wire \mexu/_0015_ ;
wire \mexu/_0016_ ;
wire \mexu/_0017_ ;
wire \mexu/_0018_ ;
wire \mexu/_0019_ ;
wire \mexu/_0020_ ;
wire \mexu/_0021_ ;
wire \mexu/_0022_ ;
wire \mexu/_0023_ ;
wire \mexu/_0024_ ;
wire \mexu/_0025_ ;
wire \mexu/_0026_ ;
wire \mexu/_0027_ ;
wire \mexu/_0028_ ;
wire \mexu/_0029_ ;
wire \mexu/_0030_ ;
wire \mexu/_0031_ ;
wire \mexu/_0032_ ;
wire \mexu/_0033_ ;
wire \mexu/_0034_ ;
wire \mexu/_0035_ ;
wire \mexu/_0036_ ;
wire \mexu/_0037_ ;
wire \mexu/_0038_ ;
wire \mexu/_0039_ ;
wire \mexu/_0040_ ;
wire \mexu/_0041_ ;
wire \mexu/_0042_ ;
wire \mexu/_0043_ ;
wire \mexu/_0044_ ;
wire \mexu/_0045_ ;
wire \mexu/_0046_ ;
wire \mexu/_0047_ ;
wire \mexu/_0048_ ;
wire \mexu/_0049_ ;
wire \mexu/_0050_ ;
wire \mexu/_0051_ ;
wire \mexu/_0052_ ;
wire \mexu/_0053_ ;
wire \mexu/_0054_ ;
wire \mexu/_0055_ ;
wire \mexu/_0056_ ;
wire \mexu/_0057_ ;
wire \mexu/_0058_ ;
wire \mexu/_0059_ ;
wire \mexu/_0060_ ;
wire \mexu/_0061_ ;
wire \mexu/_0062_ ;
wire \mexu/_0063_ ;
wire \mexu/_0064_ ;
wire \mexu/_0065_ ;
wire \mexu/_0066_ ;
wire \mexu/_0067_ ;
wire \mexu/_0068_ ;
wire \mexu/_0069_ ;
wire \mexu/_0070_ ;
wire \mexu/_0071_ ;
wire \mexu/_0072_ ;
wire \mexu/_0073_ ;
wire \mexu/_0074_ ;
wire \mexu/_0075_ ;
wire \mexu/_0076_ ;
wire \mexu/_0077_ ;
wire \mexu/_0078_ ;
wire \mexu/_0079_ ;
wire \mexu/_0080_ ;
wire \mexu/_0081_ ;
wire \mexu/_0082_ ;
wire \mexu/_0083_ ;
wire \mexu/_0084_ ;
wire \mexu/_0085_ ;
wire \mexu/_0086_ ;
wire \mexu/_0087_ ;
wire \mexu/_0088_ ;
wire \mexu/_0089_ ;
wire \mexu/_0090_ ;
wire \mexu/_0091_ ;
wire \mexu/_0092_ ;
wire \mexu/_0093_ ;
wire \mexu/_0094_ ;
wire \mexu/_0095_ ;
wire \mexu/_0096_ ;
wire \mexu/_0097_ ;
wire \mexu/_0098_ ;
wire \mexu/_0099_ ;
wire \mexu/_0100_ ;
wire \mexu/_0101_ ;
wire \mexu/_0102_ ;
wire \mexu/_0103_ ;
wire \mexu/_0104_ ;
wire \mexu/_0105_ ;
wire \mexu/_0106_ ;
wire \mexu/_0107_ ;
wire \mexu/_0108_ ;
wire \mexu/_0109_ ;
wire \mexu/_0110_ ;
wire \mexu/_0111_ ;
wire \mexu/_0112_ ;
wire \mexu/_0113_ ;
wire \mexu/_0114_ ;
wire \mexu/_0115_ ;
wire \mexu/_0116_ ;
wire \mexu/_0117_ ;
wire \mexu/_0118_ ;
wire \mexu/_0119_ ;
wire \mexu/_0120_ ;
wire \mexu/_0121_ ;
wire \mexu/_0122_ ;
wire \mexu/_0123_ ;
wire \mexu/_0124_ ;
wire \mexu/_0125_ ;
wire \mexu/_0126_ ;
wire \mexu/_0127_ ;
wire \mexu/_0128_ ;
wire \mexu/_0129_ ;
wire \mexu/_0130_ ;
wire \mexu/_0131_ ;
wire \mexu/_0132_ ;
wire \mexu/_0133_ ;
wire \mexu/_0134_ ;
wire \mexu/_0135_ ;
wire \mexu/_0136_ ;
wire \mexu/_0137_ ;
wire \mexu/_0138_ ;
wire \mexu/_0139_ ;
wire \mexu/_0140_ ;
wire \mexu/_0141_ ;
wire \mexu/_0142_ ;
wire \mexu/_0143_ ;
wire \mexu/_0144_ ;
wire \mexu/_0145_ ;
wire \mexu/_0146_ ;
wire \mexu/_0147_ ;
wire \mexu/_0148_ ;
wire \mexu/_0149_ ;
wire \mexu/_0150_ ;
wire \mexu/_0151_ ;
wire \mexu/_0152_ ;
wire \mexu/_0153_ ;
wire \mexu/_0154_ ;
wire \mexu/_0155_ ;
wire \mexu/_0156_ ;
wire \mexu/_0157_ ;
wire \mexu/_0158_ ;
wire \mexu/_0159_ ;
wire \mexu/_0160_ ;
wire \mexu/_0161_ ;
wire \mexu/_0162_ ;
wire \mexu/_0163_ ;
wire \mexu/_0164_ ;
wire \mexu/_0165_ ;
wire \mexu/_0166_ ;
wire \mexu/_0167_ ;
wire \mexu/_0168_ ;
wire \mexu/_0169_ ;
wire \mexu/_0170_ ;
wire \mexu/_0171_ ;
wire \mexu/_0172_ ;
wire \mexu/_0173_ ;
wire \mexu/_0174_ ;
wire \mexu/_0175_ ;
wire \mexu/_0176_ ;
wire \mexu/_0177_ ;
wire \mexu/_0178_ ;
wire \mexu/_0179_ ;
wire \mexu/_0180_ ;
wire \mexu/_0181_ ;
wire \mexu/_0182_ ;
wire \mexu/_0183_ ;
wire \mexu/_0184_ ;
wire \mexu/_0185_ ;
wire \mexu/_0186_ ;
wire \mexu/_0187_ ;
wire \mexu/_0188_ ;
wire \mexu/_0189_ ;
wire \mexu/_0190_ ;
wire \mexu/_0191_ ;
wire \mexu/_0192_ ;
wire \mexu/_0193_ ;
wire \mexu/_0194_ ;
wire \mexu/_0195_ ;
wire \mexu/_0196_ ;
wire \mexu/_0197_ ;
wire \mexu/_0198_ ;
wire \mexu/_0199_ ;
wire \mexu/_0200_ ;
wire \mexu/_0201_ ;
wire \mexu/_0202_ ;
wire \mexu/_0203_ ;
wire \mexu/_0204_ ;
wire \mexu/_0205_ ;
wire \mexu/_0206_ ;
wire \mexu/_0207_ ;
wire \mexu/_0208_ ;
wire \mexu/_0209_ ;
wire \mexu/_0210_ ;
wire \mexu/_0211_ ;
wire \mexu/_0212_ ;
wire \mexu/_0213_ ;
wire \mexu/_0214_ ;
wire \mexu/_0215_ ;
wire \mexu/_0216_ ;
wire \mexu/_0217_ ;
wire \mexu/_0218_ ;
wire \mexu/_0219_ ;
wire \mexu/_0220_ ;
wire \mexu/_0221_ ;
wire \mexu/_0222_ ;
wire \mexu/_0223_ ;
wire \mexu/_0224_ ;
wire \mexu/_0225_ ;
wire \mexu/_0226_ ;
wire \mexu/_0227_ ;
wire \mexu/_0228_ ;
wire \mexu/_0229_ ;
wire \mexu/_0230_ ;
wire \mexu/_0231_ ;
wire \mexu/_0232_ ;
wire \mexu/_0233_ ;
wire \mexu/_0234_ ;
wire \mexu/_0235_ ;
wire \mexu/_0236_ ;
wire \mexu/_0237_ ;
wire \mexu/_0238_ ;
wire \mexu/_0239_ ;
wire \mexu/_0240_ ;
wire \mexu/_0241_ ;
wire \mexu/_0242_ ;
wire \mexu/_0243_ ;
wire \mexu/_0244_ ;
wire \mexu/_0245_ ;
wire \mexu/_0246_ ;
wire \mexu/_0247_ ;
wire \mexu/_0248_ ;
wire \mexu/_0249_ ;
wire \mexu/_0250_ ;
wire \mexu/_0251_ ;
wire \mexu/_0252_ ;
wire \mexu/_0253_ ;
wire \mexu/_0254_ ;
wire \mexu/_0255_ ;
wire \mexu/_0256_ ;
wire \mexu/_0257_ ;
wire \mexu/_0258_ ;
wire \mexu/_0259_ ;
wire \mexu/_0260_ ;
wire \mexu/_0261_ ;
wire \mexu/_0262_ ;
wire \mexu/_0263_ ;
wire \mexu/_0264_ ;
wire \mexu/_0265_ ;
wire \mexu/_0266_ ;
wire \mexu/_0267_ ;
wire \mexu/_0268_ ;
wire \mexu/_0269_ ;
wire \mexu/_0270_ ;
wire \mexu/_0271_ ;
wire \mexu/_0272_ ;
wire \mexu/_0273_ ;
wire \mexu/_0274_ ;
wire \mexu/_0275_ ;
wire \mexu/_0276_ ;
wire \mexu/_0277_ ;
wire \mexu/_0278_ ;
wire \mexu/_0279_ ;
wire \mexu/_0280_ ;
wire \mexu/_0281_ ;
wire \mexu/_0282_ ;
wire \mexu/_0283_ ;
wire \mexu/_0284_ ;
wire \mexu/_0285_ ;
wire \mexu/_0286_ ;
wire \mexu/_0287_ ;
wire \mexu/_0288_ ;
wire \mexu/_0289_ ;
wire \mexu/_0290_ ;
wire \mexu/_0291_ ;
wire \mexu/_0292_ ;
wire \mexu/_0293_ ;
wire \mexu/_0294_ ;
wire \mexu/_0295_ ;
wire \mexu/_0296_ ;
wire \mexu/_0297_ ;
wire \mexu/_0298_ ;
wire \mexu/_0299_ ;
wire \mexu/_0300_ ;
wire \mexu/_0301_ ;
wire \mexu/_0302_ ;
wire \mexu/_0303_ ;
wire \mexu/_0304_ ;
wire \mexu/_0305_ ;
wire \mexu/_0306_ ;
wire \mexu/_0307_ ;
wire \mexu/_0308_ ;
wire \mexu/_0309_ ;
wire \mexu/_0310_ ;
wire \mexu/_0311_ ;
wire \mexu/_0312_ ;
wire \mexu/_0313_ ;
wire \mexu/_0314_ ;
wire \mexu/_0315_ ;
wire \mexu/_0316_ ;
wire \mexu/_0317_ ;
wire \mexu/_0318_ ;
wire \mexu/_0319_ ;
wire \mexu/_0320_ ;
wire \mexu/_0321_ ;
wire \mexu/_0322_ ;
wire \mexu/_0323_ ;
wire \mexu/_0324_ ;
wire \mexu/_0325_ ;
wire \mexu/_0326_ ;
wire \mexu/_0327_ ;
wire \mexu/_0328_ ;
wire \mexu/_0329_ ;
wire \mexu/_0330_ ;
wire \mexu/_0331_ ;
wire \mexu/_0332_ ;
wire \mexu/_0333_ ;
wire \mexu/_0334_ ;
wire \mexu/_0335_ ;
wire \mexu/_0336_ ;
wire \mexu/_0337_ ;
wire \mexu/_0338_ ;
wire \mexu/_0339_ ;
wire \mexu/_0340_ ;
wire \mexu/_0341_ ;
wire \mexu/_0342_ ;
wire \mexu/_0343_ ;
wire \mexu/_0344_ ;
wire \mexu/_0345_ ;
wire \mexu/_0346_ ;
wire \mexu/_0347_ ;
wire \mexu/_0348_ ;
wire \mexu/_0349_ ;
wire \mexu/_0350_ ;
wire \mexu/_0351_ ;
wire \mexu/_0352_ ;
wire \mexu/_0353_ ;
wire \mexu/_0354_ ;
wire \mexu/_0355_ ;
wire \mexu/_0356_ ;
wire \mexu/_0357_ ;
wire \mexu/_0358_ ;
wire \mexu/_0359_ ;
wire \mexu/_0360_ ;
wire \mexu/_0361_ ;
wire \mexu/_0362_ ;
wire \mexu/_0363_ ;
wire \mexu/_0364_ ;
wire \mexu/_0365_ ;
wire \mexu/_0366_ ;
wire \mexu/_0367_ ;
wire \mexu/_0368_ ;
wire \mexu/_0369_ ;
wire \mexu/_0370_ ;
wire \mexu/_0371_ ;
wire \mexu/_0372_ ;
wire \mexu/_0373_ ;
wire \mexu/_0374_ ;
wire \mexu/_0375_ ;
wire \mexu/_0376_ ;
wire \mexu/_0377_ ;
wire \mexu/_0378_ ;
wire \mexu/_0379_ ;
wire \mexu/_0380_ ;
wire \mexu/_0381_ ;
wire \mexu/_0382_ ;
wire \mexu/_0383_ ;
wire \mexu/_0384_ ;
wire \mexu/_0385_ ;
wire \mexu/_0386_ ;
wire \mexu/_0387_ ;
wire \mexu/_0388_ ;
wire \mexu/_0389_ ;
wire \mexu/_0390_ ;
wire \mexu/_0391_ ;
wire \mexu/_0392_ ;
wire \mexu/_0393_ ;
wire \mexu/_0394_ ;
wire \mexu/_0395_ ;
wire \mexu/_0396_ ;
wire \mexu/_0397_ ;
wire \mexu/_0398_ ;
wire \mexu/_0399_ ;
wire \mexu/_0400_ ;
wire \mexu/_0401_ ;
wire \mexu/_0402_ ;
wire \mexu/_0403_ ;
wire \mexu/_0404_ ;
wire \mexu/_0405_ ;
wire \mexu/_0406_ ;
wire \mexu/_0407_ ;
wire \mexu/_0408_ ;
wire \mexu/_0409_ ;
wire \mexu/_0410_ ;
wire \mexu/_0411_ ;
wire \mexu/_0412_ ;
wire \mexu/_0413_ ;
wire \mexu/_0414_ ;
wire \mexu/_0415_ ;
wire \mexu/_0416_ ;
wire \mexu/_0417_ ;
wire \mexu/_0418_ ;
wire \mexu/_0419_ ;
wire \mexu/_0420_ ;
wire \mexu/_0421_ ;
wire \mexu/_0422_ ;
wire \mexu/_0423_ ;
wire \mexu/_0424_ ;
wire \mexu/_0425_ ;
wire \mexu/_0426_ ;
wire \mexu/_0427_ ;
wire \mexu/_0428_ ;
wire \mexu/_0429_ ;
wire \mexu/_0430_ ;
wire \mexu/_0431_ ;
wire \mexu/_0432_ ;
wire \mexu/_0433_ ;
wire \mexu/_0434_ ;
wire \mexu/_0435_ ;
wire \mexu/_0436_ ;
wire \mexu/_0437_ ;
wire \mexu/_0438_ ;
wire \mexu/_0439_ ;
wire \mexu/_0440_ ;
wire \mexu/_0441_ ;
wire \mexu/_0442_ ;
wire \mexu/_0443_ ;
wire \mexu/_0444_ ;
wire \mexu/_0445_ ;
wire \mexu/_0446_ ;
wire \mexu/_0447_ ;
wire \mexu/_0448_ ;
wire \mexu/_0449_ ;
wire \mexu/_0450_ ;
wire \mexu/_0451_ ;
wire \mexu/_0452_ ;
wire \mexu/_0453_ ;
wire \mexu/_0454_ ;
wire \mexu/_0455_ ;
wire \mexu/_0456_ ;
wire \mexu/_0457_ ;
wire \mexu/_0458_ ;
wire \mexu/_0459_ ;
wire \mexu/_0460_ ;
wire \mexu/_0461_ ;
wire \mexu/_0462_ ;
wire \mexu/_0463_ ;
wire \mexu/_0464_ ;
wire \mexu/_0465_ ;
wire \mexu/_0466_ ;
wire \mexu/_0467_ ;
wire \mexu/_0468_ ;
wire \mexu/_0469_ ;
wire \mexu/_0470_ ;
wire \mexu/_0471_ ;
wire \mexu/_0472_ ;
wire \mexu/_0473_ ;
wire \mexu/_0474_ ;
wire \mexu/_0475_ ;
wire \mexu/_0476_ ;
wire \mexu/_0477_ ;
wire \mexu/_0478_ ;
wire \mexu/_0479_ ;
wire \mexu/_0480_ ;
wire \mexu/_0481_ ;
wire \mexu/_0482_ ;
wire \mexu/_0483_ ;
wire \mexu/_0484_ ;
wire \mexu/_0485_ ;
wire \mexu/_0486_ ;
wire \mexu/_0487_ ;
wire \mexu/_0488_ ;
wire \mexu/_0489_ ;
wire \mexu/_0490_ ;
wire \mexu/_0491_ ;
wire \mexu/_0492_ ;
wire \mexu/_0493_ ;
wire \mexu/_0494_ ;
wire \mexu/_0495_ ;
wire \mexu/_0496_ ;
wire \mexu/_0497_ ;
wire \mexu/_0498_ ;
wire \mexu/_0499_ ;
wire \mexu/_0500_ ;
wire \mexu/_0501_ ;
wire \mexu/_0502_ ;
wire \mexu/_0503_ ;
wire \mexu/_0504_ ;
wire \mexu/_0505_ ;
wire \mexu/_0506_ ;
wire \mexu/_0507_ ;
wire \mexu/_0508_ ;
wire \mexu/_0509_ ;
wire \mexu/_0510_ ;
wire \mexu/_0511_ ;
wire \mexu/_0512_ ;
wire \mexu/_0513_ ;
wire \mexu/_0514_ ;
wire \mexu/_0515_ ;
wire \mexu/_0516_ ;
wire \mexu/_0517_ ;
wire \mexu/_0518_ ;
wire \mexu/_0519_ ;
wire \mexu/_0520_ ;
wire \mexu/_0521_ ;
wire \mexu/_0522_ ;
wire \mexu/_0523_ ;
wire \mexu/_0524_ ;
wire \mexu/_0525_ ;
wire \mexu/_0526_ ;
wire \mexu/_0527_ ;
wire \mexu/_0528_ ;
wire \mexu/_0529_ ;
wire \mexu/_0530_ ;
wire \mexu/_0531_ ;
wire \mexu/_0532_ ;
wire \mexu/_0533_ ;
wire \mexu/_0534_ ;
wire \mexu/_0535_ ;
wire \mexu/_0536_ ;
wire \mexu/_0537_ ;
wire \mexu/_0538_ ;
wire \mexu/_0539_ ;
wire \mexu/_0540_ ;
wire \mexu/_0541_ ;
wire \mexu/_0542_ ;
wire \mexu/_0543_ ;
wire \mexu/_0544_ ;
wire \mexu/_0545_ ;
wire \mexu/_0546_ ;
wire \mexu/_0547_ ;
wire \mexu/_0548_ ;
wire \mexu/_0549_ ;
wire \mexu/_0550_ ;
wire \mexu/_0551_ ;
wire \mexu/_0552_ ;
wire \mexu/_0553_ ;
wire \mexu/_0554_ ;
wire \mexu/_0555_ ;
wire \mexu/_0556_ ;
wire \mexu/_0557_ ;
wire \mexu/_0558_ ;
wire \mexu/_0559_ ;
wire \mexu/_0560_ ;
wire \mexu/_0561_ ;
wire \mexu/_0562_ ;
wire \mexu/_0563_ ;
wire \mexu/_0564_ ;
wire \mexu/_0565_ ;
wire \mexu/_0566_ ;
wire \mexu/_0567_ ;
wire \mexu/_0568_ ;
wire \mexu/_0569_ ;
wire \mexu/_0570_ ;
wire \mexu/_0571_ ;
wire \mexu/_0572_ ;
wire \mexu/_0573_ ;
wire \mexu/_0574_ ;
wire \mexu/_0575_ ;
wire \mexu/_0576_ ;
wire \mexu/_0577_ ;
wire \mexu/_0578_ ;
wire \mexu/_0579_ ;
wire \mexu/_0580_ ;
wire \mexu/_0581_ ;
wire \mexu/_0582_ ;
wire \mexu/_0583_ ;
wire \mexu/_0584_ ;
wire \mexu/_0585_ ;
wire \mexu/_0586_ ;
wire \mexu/_0587_ ;
wire \mexu/_0588_ ;
wire \mexu/_0589_ ;
wire \mexu/_0590_ ;
wire \mexu/_0591_ ;
wire \mexu/_0592_ ;
wire \mexu/_0593_ ;
wire \mexu/_0594_ ;
wire \mexu/_0595_ ;
wire \mexu/_0596_ ;
wire \mexu/_0597_ ;
wire \mexu/_0598_ ;
wire \mexu/_0599_ ;
wire \mexu/_0600_ ;
wire \mexu/_0601_ ;
wire \mexu/_0602_ ;
wire \mexu/_0603_ ;
wire \mexu/_0604_ ;
wire \mexu/_0605_ ;
wire \mexu/_0606_ ;
wire \mexu/_0607_ ;
wire \mexu/_0608_ ;
wire \mexu/_0609_ ;
wire \mexu/_0610_ ;
wire \mexu/_0611_ ;
wire \mexu/_0612_ ;
wire \mexu/_0613_ ;
wire \mexu/_0614_ ;
wire \mexu/_0615_ ;
wire \mexu/_0616_ ;
wire \mexu/_0617_ ;
wire \mexu/_0618_ ;
wire \mexu/_0619_ ;
wire \mexu/_0620_ ;
wire \mexu/_0621_ ;
wire \mexu/_0622_ ;
wire \mexu/_0623_ ;
wire \mexu/_0624_ ;
wire \mexu/_0625_ ;
wire \mexu/_0626_ ;
wire \mexu/_0627_ ;
wire \mexu/_0628_ ;
wire \mexu/_0629_ ;
wire \mexu/_0630_ ;
wire \mexu/_0631_ ;
wire \mexu/_0632_ ;
wire \mexu/_0633_ ;
wire \mexu/_0634_ ;
wire \mexu/_0635_ ;
wire \mexu/_0636_ ;
wire \mexu/_0637_ ;
wire \mexu/_0638_ ;
wire \mexu/_0639_ ;
wire \mexu/_0640_ ;
wire \mexu/_0641_ ;
wire \mexu/_0642_ ;
wire \mexu/_0643_ ;
wire \mexu/_0644_ ;
wire \mexu/_0645_ ;
wire \mexu/_0646_ ;
wire \mexu/_0647_ ;
wire \mexu/_0648_ ;
wire \mexu/_0649_ ;
wire \mexu/_0650_ ;
wire \mexu/_0651_ ;
wire \mexu/_0652_ ;
wire \mexu/_0653_ ;
wire \mexu/_0654_ ;
wire \mexu/_0655_ ;
wire \mexu/_0656_ ;
wire \mexu/_0657_ ;
wire \mexu/_0658_ ;
wire \mexu/_0659_ ;
wire \mexu/_0660_ ;
wire \mexu/_0661_ ;
wire \mexu/_0662_ ;
wire \mexu/_0663_ ;
wire \mexu/_0664_ ;
wire \mexu/_0665_ ;
wire \mexu/_0666_ ;
wire \mexu/_0667_ ;
wire \mexu/_0668_ ;
wire \mexu/_0669_ ;
wire \mexu/_0670_ ;
wire \mexu/_0671_ ;
wire \mexu/_0672_ ;
wire \mexu/_0673_ ;
wire \mexu/_0674_ ;
wire \mexu/_0675_ ;
wire \mexu/_0676_ ;
wire \mexu/_0677_ ;
wire \mexu/_0678_ ;
wire \mexu/_0679_ ;
wire \mexu/_0680_ ;
wire \mexu/_0681_ ;
wire \mexu/_0682_ ;
wire \mexu/_0683_ ;
wire \mexu/_0684_ ;
wire \mexu/_0685_ ;
wire \mexu/_0686_ ;
wire \mexu/_0687_ ;
wire \mexu/_0688_ ;
wire \mexu/_0689_ ;
wire \mexu/_0690_ ;
wire \mexu/_0691_ ;
wire \mexu/_0692_ ;
wire \mexu/_0693_ ;
wire \mexu/_0694_ ;
wire \mexu/_0695_ ;
wire \mexu/_0696_ ;
wire \mexu/_0697_ ;
wire \mexu/_0698_ ;
wire \mexu/_0699_ ;
wire \mexu/_0700_ ;
wire \mexu/_0701_ ;
wire \mexu/_0702_ ;
wire \mexu/_0703_ ;
wire \mexu/_0704_ ;
wire \mexu/_0705_ ;
wire \mexu/_0706_ ;
wire \mexu/_0707_ ;
wire \mexu/_0708_ ;
wire \mexu/_0709_ ;
wire \mexu/_0710_ ;
wire \mexu/_0711_ ;
wire \mexu/_0712_ ;
wire \mexu/_0713_ ;
wire \mexu/_0714_ ;
wire \mexu/_0715_ ;
wire \mexu/_0716_ ;
wire \mexu/_0717_ ;
wire \mexu/_0718_ ;
wire \mexu/_0719_ ;
wire \mexu/_0720_ ;
wire \mexu/_0721_ ;
wire \mexu/_0722_ ;
wire \mexu/_0723_ ;
wire \mexu/_0724_ ;
wire \mexu/_0725_ ;
wire \mexu/_0726_ ;
wire \mexu/_0727_ ;
wire \mexu/_0728_ ;
wire \mexu/_0729_ ;
wire \mexu/_0730_ ;
wire \mexu/_0731_ ;
wire \mexu/_0732_ ;
wire \mexu/_0733_ ;
wire \mexu/_0734_ ;
wire \mexu/_0735_ ;
wire \mexu/_0736_ ;
wire \mexu/_0737_ ;
wire \mexu/_0738_ ;
wire \mexu/_0739_ ;
wire \mexu/_0740_ ;
wire \mexu/_0741_ ;
wire \mexu/_0742_ ;
wire \mexu/_0743_ ;
wire \mexu/_0744_ ;
wire \mexu/_0745_ ;
wire \mexu/_0746_ ;
wire \mexu/_0747_ ;
wire \mexu/_0748_ ;
wire \mexu/_0749_ ;
wire \mexu/_0750_ ;
wire \mexu/_0751_ ;
wire \mexu/_0752_ ;
wire \mexu/_0753_ ;
wire \mexu/_0754_ ;
wire \mexu/_0755_ ;
wire \mexu/_0756_ ;
wire \mexu/_0757_ ;
wire \mexu/_0758_ ;
wire \mexu/_0759_ ;
wire \mexu/_0760_ ;
wire \mexu/_0761_ ;
wire \mexu/_0762_ ;
wire \mexu/_0763_ ;
wire \mexu/_0764_ ;
wire \mexu/_0765_ ;
wire \mexu/_0766_ ;
wire \mexu/_0767_ ;
wire \mexu/_0768_ ;
wire \mexu/_0769_ ;
wire \mexu/_0770_ ;
wire \mexu/_0771_ ;
wire \mexu/_0772_ ;
wire \mexu/_0773_ ;
wire \mexu/_0774_ ;
wire \mexu/_0775_ ;
wire \mexu/_0776_ ;
wire \mexu/_0777_ ;
wire \mexu/_0778_ ;
wire \mexu/_0779_ ;
wire \mexu/_0780_ ;
wire \mexu/_0781_ ;
wire \mexu/_0782_ ;
wire \mexu/_0783_ ;
wire \mexu/_0784_ ;
wire \mexu/_0785_ ;
wire \mexu/_0786_ ;
wire \mexu/_0787_ ;
wire \mexu/_0788_ ;
wire \mexu/_0789_ ;
wire \mexu/_0790_ ;
wire \mexu/_0791_ ;
wire \mexu/_0792_ ;
wire \mexu/_0793_ ;
wire \mexu/_0794_ ;
wire \mexu/_0795_ ;
wire \mexu/_0796_ ;
wire \mexu/_0797_ ;
wire \mexu/_0798_ ;
wire \mexu/_0799_ ;
wire \mexu/_0800_ ;
wire \mexu/_0801_ ;
wire \mexu/_0802_ ;
wire \mexu/_0803_ ;
wire \mexu/_0804_ ;
wire \mexu/_0805_ ;
wire \mexu/_0806_ ;
wire \mexu/_0807_ ;
wire \mexu/_0808_ ;
wire \mexu/_0809_ ;
wire \mexu/_0810_ ;
wire \mexu/_0811_ ;
wire \mexu/_0812_ ;
wire \mexu/_0813_ ;
wire \mexu/_0814_ ;
wire \mexu/_0815_ ;
wire \mexu/_0816_ ;
wire \mexu/_0817_ ;
wire \mexu/_0818_ ;
wire \mexu/_0819_ ;
wire \mexu/_0820_ ;
wire \mexu/_0821_ ;
wire \mexu/_0822_ ;
wire \mexu/_0823_ ;
wire \mexu/_0824_ ;
wire \mexu/_0825_ ;
wire \mexu/_0826_ ;
wire \mexu/_0827_ ;
wire \mexu/_0828_ ;
wire \mexu/_0829_ ;
wire \mexu/_0830_ ;
wire \mexu/_0831_ ;
wire \mexu/_0832_ ;
wire \mexu/_0833_ ;
wire \mexu/_0834_ ;
wire \mexu/_0835_ ;
wire \mexu/_0836_ ;
wire \mexu/_0837_ ;
wire \mexu/_0838_ ;
wire \mexu/_0839_ ;
wire \mexu/_0840_ ;
wire \mexu/_0841_ ;
wire \mexu/_0842_ ;
wire \mexu/_0843_ ;
wire \mexu/_0844_ ;
wire \mexu/_0845_ ;
wire \mexu/_0846_ ;
wire \mexu/_0847_ ;
wire \mexu/_0848_ ;
wire \mexu/_0849_ ;
wire \mexu/_0850_ ;
wire \mexu/_0851_ ;
wire \mexu/_0852_ ;
wire \mexu/_0853_ ;
wire \mexu/_0854_ ;
wire \mexu/_0855_ ;
wire \mexu/_0856_ ;
wire \mexu/_0857_ ;
wire \mexu/_0858_ ;
wire \mexu/_0859_ ;
wire \mexu/_0860_ ;
wire \mexu/_0861_ ;
wire \mexu/_0862_ ;
wire \mexu/_0863_ ;
wire \mexu/_0864_ ;
wire \mexu/_0865_ ;
wire \mexu/_0866_ ;
wire \mexu/_0867_ ;
wire \mexu/_0868_ ;
wire \mexu/_0869_ ;
wire \mexu/_0870_ ;
wire \mexu/_0871_ ;
wire \mexu/_0872_ ;
wire \mexu/_0873_ ;
wire \mexu/_0874_ ;
wire \mexu/_0875_ ;
wire \mexu/_0876_ ;
wire \mexu/_0877_ ;
wire \mexu/_0878_ ;
wire \mexu/_0879_ ;
wire \mexu/_0880_ ;
wire \mexu/_0881_ ;
wire \mexu/_0882_ ;
wire \mexu/_0883_ ;
wire \mexu/_0884_ ;
wire \mexu/_0885_ ;
wire \mexu/_0886_ ;
wire \mexu/_0887_ ;
wire \mexu/_0888_ ;
wire \mexu/_0889_ ;
wire \mexu/_0890_ ;
wire \mexu/_0891_ ;
wire \mexu/_0892_ ;
wire \mexu/_0893_ ;
wire \mexu/_0894_ ;
wire \mexu/_0895_ ;
wire \mexu/_0896_ ;
wire \mexu/_0897_ ;
wire \mexu/_0898_ ;
wire \mexu/_0899_ ;
wire \mexu/_0900_ ;
wire \mexu/_0901_ ;
wire \mexu/_0902_ ;
wire \mexu/_0903_ ;
wire \mexu/_0904_ ;
wire \mexu/_0905_ ;
wire \mexu/_0906_ ;
wire \mexu/_0907_ ;
wire \mexu/_0908_ ;
wire \mexu/_0909_ ;
wire \mexu/_0910_ ;
wire \mexu/_0911_ ;
wire \mexu/_0912_ ;
wire \mexu/_0913_ ;
wire \mexu/_0914_ ;
wire \mexu/_0915_ ;
wire \mexu/_0916_ ;
wire \mexu/_0917_ ;
wire \mexu/_0918_ ;
wire \mexu/_0919_ ;
wire \mexu/_0920_ ;
wire \mexu/_0921_ ;
wire \mexu/_0922_ ;
wire \mexu/_0923_ ;
wire \mexu/_0924_ ;
wire \mexu/_0925_ ;
wire \mexu/_0926_ ;
wire \mexu/_0927_ ;
wire \mexu/_0928_ ;
wire \mexu/_0929_ ;
wire \mexu/_0930_ ;
wire \mexu/_0931_ ;
wire \mexu/_0932_ ;
wire \mexu/_0933_ ;
wire \mexu/_0934_ ;
wire \mexu/_0935_ ;
wire \mexu/_0936_ ;
wire \mexu/_0937_ ;
wire \mexu/_0938_ ;
wire \mexu/_0939_ ;
wire \mexu/_0940_ ;
wire \mexu/_0941_ ;
wire \mexu/_0942_ ;
wire \mexu/_0943_ ;
wire \mexu/_0944_ ;
wire \mexu/_0945_ ;
wire \mexu/_0946_ ;
wire \mexu/_0947_ ;
wire \mexu/_0948_ ;
wire \mexu/_0949_ ;
wire \mexu/_0950_ ;
wire \mexu/_0951_ ;
wire \mexu/_0952_ ;
wire \mexu/_0953_ ;
wire \mexu/_0954_ ;
wire \mexu/_0955_ ;
wire \mexu/_0956_ ;
wire \mexu/_0957_ ;
wire \mexu/_0958_ ;
wire \mexu/_0959_ ;
wire \mexu/_0960_ ;
wire \mexu/_0961_ ;
wire \mexu/_0962_ ;
wire \mexu/_0963_ ;
wire \mexu/_0964_ ;
wire \mexu/_0965_ ;
wire \mexu/_0966_ ;
wire \mexu/_0967_ ;
wire \mexu/_0968_ ;
wire \mexu/_0969_ ;
wire \mexu/_0970_ ;
wire \mexu/_0971_ ;
wire \mexu/_0972_ ;
wire \mexu/_0973_ ;
wire \mexu/_0974_ ;
wire \mexu/_0975_ ;
wire \mexu/_0976_ ;
wire \mexu/_0977_ ;
wire \mexu/_0978_ ;
wire \mexu/_0979_ ;
wire \mexu/_0980_ ;
wire \mexu/_0981_ ;
wire \mexu/_0982_ ;
wire \mexu/_0983_ ;
wire \mexu/_0984_ ;
wire \mexu/_0985_ ;
wire \mexu/_0986_ ;
wire \mexu/_0987_ ;
wire \mexu/_0988_ ;
wire \mexu/_0989_ ;
wire \mexu/_0990_ ;
wire \mexu/_0991_ ;
wire \mexu/_0992_ ;
wire \mexu/_0993_ ;
wire \mexu/_0994_ ;
wire \mexu/_0995_ ;
wire \mexu/_0996_ ;
wire \mexu/_0997_ ;
wire \mexu/_0998_ ;
wire \mexu/_0999_ ;
wire \mexu/_1000_ ;
wire \mexu/_1001_ ;
wire \mexu/_1002_ ;
wire \mexu/_1003_ ;
wire \mexu/_1004_ ;
wire \mexu/_1005_ ;
wire \mexu/_1006_ ;
wire \mexu/_1007_ ;
wire \mexu/_1008_ ;
wire \mexu/_1009_ ;
wire \mexu/_1010_ ;
wire \mexu/_1011_ ;
wire \mexu/_1012_ ;
wire \mexu/_1013_ ;
wire \mexu/_1014_ ;
wire \mexu/_1015_ ;
wire \mexu/_1016_ ;
wire \mexu/_1017_ ;
wire \mexu/_1018_ ;
wire \mexu/_1019_ ;
wire \mexu/_1020_ ;
wire \mexu/_1021_ ;
wire \mexu/_1022_ ;
wire \mexu/_1023_ ;
wire \mexu/_1024_ ;
wire \mexu/_1025_ ;
wire \mexu/_1026_ ;
wire \mexu/_1027_ ;
wire \mexu/_1028_ ;
wire \mexu/_1029_ ;
wire \mexu/_1030_ ;
wire \mexu/_1031_ ;
wire \mexu/_1032_ ;
wire \mexu/_1033_ ;
wire \mexu/_1034_ ;
wire \mexu/_1035_ ;
wire \mexu/_1036_ ;
wire \mexu/_1037_ ;
wire \mexu/_1038_ ;
wire \mexu/_1039_ ;
wire \mexu/_1040_ ;
wire \mexu/_1041_ ;
wire \mexu/_1042_ ;
wire \mexu/_1043_ ;
wire \mexu/_1044_ ;
wire \mexu/_1045_ ;
wire \mexu/_1046_ ;
wire \mexu/_1047_ ;
wire \mexu/_1048_ ;
wire \mexu/_1049_ ;
wire \mexu/_1050_ ;
wire \mexu/_1051_ ;
wire \mexu/_1052_ ;
wire \mexu/_1053_ ;
wire \mexu/_1054_ ;
wire \mexu/_1055_ ;
wire \mexu/_1056_ ;
wire \mexu/_1057_ ;
wire \mexu/_1058_ ;
wire \mexu/_1059_ ;
wire \mexu/_1060_ ;
wire \mexu/_1061_ ;
wire \mexu/_1062_ ;
wire \mexu/_1063_ ;
wire \mexu/_1064_ ;
wire \mexu/_1065_ ;
wire \mexu/_1066_ ;
wire \mexu/_1067_ ;
wire \mexu/_1068_ ;
wire \mexu/_1069_ ;
wire \mexu/_1070_ ;
wire \mexu/_1071_ ;
wire \mexu/_1072_ ;
wire \mexu/_1073_ ;
wire \mexu/_1074_ ;
wire \mexu/_1075_ ;
wire \mexu/_1076_ ;
wire \mexu/_1077_ ;
wire \mexu/_1078_ ;
wire \mexu/_1079_ ;
wire \mexu/_1080_ ;
wire \mexu/_1081_ ;
wire \mexu/_1082_ ;
wire \mexu/_1083_ ;
wire \mexu/_1084_ ;
wire \mexu/_1085_ ;
wire \mexu/_1086_ ;
wire \mexu/_1087_ ;
wire \mexu/_1088_ ;
wire \mexu/_1089_ ;
wire \mexu/_1090_ ;
wire \mexu/_1091_ ;
wire \mexu/_1092_ ;
wire \mexu/_1093_ ;
wire \midu/_000_ ;
wire \midu/_001_ ;
wire \midu/_002_ ;
wire \midu/_003_ ;
wire \midu/_004_ ;
wire \midu/_005_ ;
wire \midu/_006_ ;
wire \midu/_007_ ;
wire \midu/_008_ ;
wire \midu/_009_ ;
wire \midu/_010_ ;
wire \midu/_011_ ;
wire \midu/_012_ ;
wire \midu/_013_ ;
wire \midu/_014_ ;
wire \midu/_015_ ;
wire \midu/_016_ ;
wire \midu/_017_ ;
wire \midu/_018_ ;
wire \midu/_019_ ;
wire \midu/_020_ ;
wire \midu/_021_ ;
wire \midu/_022_ ;
wire \midu/_023_ ;
wire \midu/_024_ ;
wire \midu/_025_ ;
wire \midu/_026_ ;
wire \midu/_027_ ;
wire \midu/_028_ ;
wire \midu/_029_ ;
wire \midu/_030_ ;
wire \midu/_031_ ;
wire \midu/_032_ ;
wire \midu/_033_ ;
wire \midu/_034_ ;
wire \midu/_035_ ;
wire \midu/_036_ ;
wire \midu/_037_ ;
wire \midu/_038_ ;
wire \midu/_039_ ;
wire \midu/_040_ ;
wire \midu/_041_ ;
wire \midu/_042_ ;
wire \midu/_043_ ;
wire \midu/_044_ ;
wire \midu/_045_ ;
wire \midu/_046_ ;
wire \midu/_047_ ;
wire \midu/_048_ ;
wire \midu/_049_ ;
wire \midu/_050_ ;
wire \midu/_051_ ;
wire \midu/_052_ ;
wire \midu/_053_ ;
wire \midu/_054_ ;
wire \midu/_055_ ;
wire \midu/_056_ ;
wire \midu/_057_ ;
wire \midu/_058_ ;
wire \midu/_059_ ;
wire \midu/_060_ ;
wire \midu/_061_ ;
wire \midu/_062_ ;
wire \midu/_063_ ;
wire \midu/_064_ ;
wire \midu/_065_ ;
wire \midu/_066_ ;
wire \midu/_067_ ;
wire \midu/_068_ ;
wire \midu/_069_ ;
wire \midu/_070_ ;
wire \midu/_071_ ;
wire \midu/_072_ ;
wire \midu/_073_ ;
wire \midu/_074_ ;
wire \midu/_075_ ;
wire \midu/_076_ ;
wire \midu/_077_ ;
wire \midu/_078_ ;
wire \midu/_079_ ;
wire \midu/_080_ ;
wire \midu/_081_ ;
wire \midu/_082_ ;
wire \midu/_083_ ;
wire \midu/_084_ ;
wire \midu/_085_ ;
wire \midu/_086_ ;
wire \midu/_087_ ;
wire \midu/_088_ ;
wire \midu/_089_ ;
wire \midu/_090_ ;
wire \midu/_091_ ;
wire \midu/_092_ ;
wire \midu/_093_ ;
wire \midu/_094_ ;
wire \midu/_095_ ;
wire \midu/_096_ ;
wire \midu/_097_ ;
wire \midu/_098_ ;
wire \midu/_099_ ;
wire \midu/_100_ ;
wire \midu/_101_ ;
wire \midu/_102_ ;
wire \midu/_103_ ;
wire \midu/_104_ ;
wire \midu/_105_ ;
wire \midu/_106_ ;
wire \midu/_107_ ;
wire \midu/_108_ ;
wire \midu/_109_ ;
wire \midu/_110_ ;
wire \midu/_111_ ;
wire \midu/_112_ ;
wire \midu/_113_ ;
wire \midu/_114_ ;
wire \midu/_115_ ;
wire \midu/_116_ ;
wire \midu/_117_ ;
wire \midu/_118_ ;
wire \midu/_119_ ;
wire \midu/_120_ ;
wire \midu/_121_ ;
wire \midu/_122_ ;
wire \midu/_123_ ;
wire \midu/_124_ ;
wire \midu/_125_ ;
wire \midu/_126_ ;
wire \midu/_127_ ;
wire \midu/_128_ ;
wire \midu/_129_ ;
wire \midu/_130_ ;
wire \mifu/_000_ ;
wire \mifu/_001_ ;
wire \mifu/_002_ ;
wire \mifu/_003_ ;
wire \mifu/_004_ ;
wire \mifu/_005_ ;
wire \mifu/_006_ ;
wire \mifu/_007_ ;
wire \mifu/_008_ ;
wire \mifu/_009_ ;
wire \mifu/_010_ ;
wire \mifu/_011_ ;
wire \mifu/_012_ ;
wire \mifu/_013_ ;
wire \mifu/_014_ ;
wire \mifu/_015_ ;
wire \mifu/_016_ ;
wire \mifu/_017_ ;
wire \mifu/_018_ ;
wire \mifu/_019_ ;
wire \mifu/_020_ ;
wire \mifu/_021_ ;
wire \mifu/_022_ ;
wire \mifu/_023_ ;
wire \mifu/_024_ ;
wire \mifu/_025_ ;
wire \mifu/_026_ ;
wire \mifu/_027_ ;
wire \mifu/_028_ ;
wire \mifu/_029_ ;
wire \mifu/_030_ ;
wire \mifu/_031_ ;
wire \mifu/_032_ ;
wire \mifu/_033_ ;
wire \mifu/_034_ ;
wire \mifu/_035_ ;
wire \mifu/_036_ ;
wire \mifu/_037_ ;
wire \mifu/_038_ ;
wire \mifu/_039_ ;
wire \mifu/_040_ ;
wire \mifu/_041_ ;
wire \mifu/_042_ ;
wire \mifu/_043_ ;
wire \mifu/_044_ ;
wire \mifu/_045_ ;
wire \mifu/_046_ ;
wire \mifu/_047_ ;
wire \mifu/_048_ ;
wire \mifu/_049_ ;
wire \mifu/_050_ ;
wire \mifu/_051_ ;
wire \mifu/_052_ ;
wire \mifu/_053_ ;
wire \mifu/_054_ ;
wire \mifu/_055_ ;
wire \mifu/_056_ ;
wire \mifu/_057_ ;
wire \mifu/_058_ ;
wire \mifu/_059_ ;
wire \mifu/_060_ ;
wire \mifu/_061_ ;
wire \mifu/_062_ ;
wire \mifu/_063_ ;
wire \mifu/_064_ ;
wire \mifu/_065_ ;
wire \mifu/_066_ ;
wire \mifu/_067_ ;
wire \mifu/_068_ ;
wire \mifu/_069_ ;
wire \mifu/_070_ ;
wire \mifu/_071_ ;
wire \mifu/_072_ ;
wire \mifu/_073_ ;
wire \mifu/_074_ ;
wire \mifu/_075_ ;
wire \mifu/_076_ ;
wire \mifu/_077_ ;
wire \mifu/_078_ ;
wire \mifu/_079_ ;
wire \mifu/_080_ ;
wire \mifu/_081_ ;
wire \mifu/_082_ ;
wire \mifu/_083_ ;
wire \mifu/_084_ ;
wire \mifu/_085_ ;
wire \mifu/_086_ ;
wire \mifu/_087_ ;
wire \mifu/_088_ ;
wire \mifu/_089_ ;
wire \mifu/_090_ ;
wire \mifu/_091_ ;
wire \mifu/_092_ ;
wire \mifu/_093_ ;
wire \mifu/_094_ ;
wire \mifu/_095_ ;
wire \mifu/_096_ ;
wire \mifu/_097_ ;
wire \mifu/_098_ ;
wire \mifu/_099_ ;
wire \mifu/_100_ ;
wire \mifu/_101_ ;
wire \mifu/_102_ ;
wire \mifu/_103_ ;
wire \mifu/_104_ ;
wire \mifu/_105_ ;
wire \mifu/_106_ ;
wire \mifu/_107_ ;
wire \mifu/_108_ ;
wire \mifu/_109_ ;
wire \mifu/_110_ ;
wire \mifu/_111_ ;
wire \mifu/_112_ ;
wire \mifu/_113_ ;
wire \mifu/_114_ ;
wire \mifu/_115_ ;
wire \mifu/_116_ ;
wire \mifu/_117_ ;
wire \mifu/_118_ ;
wire \mifu/_119_ ;
wire \mifu/_120_ ;
wire \mifu/_121_ ;
wire \mifu/_122_ ;
wire \mifu/_123_ ;
wire \mifu/_124_ ;
wire \mifu/_125_ ;
wire \mifu/_126_ ;
wire \mifu/_127_ ;
wire \mifu/_128_ ;
wire \mifu/_129_ ;
wire \mifu/_130_ ;
wire \mifu/_131_ ;
wire \mifu/_132_ ;
wire \mifu/_133_ ;
wire \mifu/_134_ ;
wire \mifu/_135_ ;
wire \mifu/_136_ ;
wire \mifu/_137_ ;
wire \mifu/_138_ ;
wire \mifu/_139_ ;
wire \mifu/_140_ ;
wire \mifu/_141_ ;
wire \mifu/_142_ ;
wire \mifu/_143_ ;
wire \mifu/_144_ ;
wire \mifu/_145_ ;
wire \mifu/_146_ ;
wire \mifu/_147_ ;
wire \mifu/_148_ ;
wire \mifu/_149_ ;
wire \mifu/_150_ ;
wire \mifu/_151_ ;
wire \mifu/_152_ ;
wire \mifu/_153_ ;
wire \mifu/_154_ ;
wire \mifu/_155_ ;
wire \mifu/_156_ ;
wire \mifu/_157_ ;
wire \mifu/_158_ ;
wire \mifu/_159_ ;
wire \mifu/_160_ ;
wire \mifu/_161_ ;
wire \mifu/_162_ ;
wire \mifu/_163_ ;
wire \mifu/_164_ ;
wire \mifu/_165_ ;
wire \mifu/_166_ ;
wire \mifu/_167_ ;
wire \mifu/_168_ ;
wire \mifu/_169_ ;
wire \mifu/_170_ ;
wire \mifu/_171_ ;
wire \mifu/_172_ ;
wire \mifu/_173_ ;
wire \mifu/_174_ ;
wire \mifu/_175_ ;
wire \mifu/_176_ ;
wire \mifu/_177_ ;
wire \mifu/_178_ ;
wire \mifu/_179_ ;
wire \mifu/_180_ ;
wire \mifu/_181_ ;
wire \mifu/_182_ ;
wire \mifu/_183_ ;
wire \mifu/_184_ ;
wire \mifu/_185_ ;
wire \mifu/_186_ ;
wire \mifu/_187_ ;
wire \mifu/_188_ ;
wire \mifu/_189_ ;
wire \mifu/_190_ ;
wire \mifu/_191_ ;
wire \mifu/_192_ ;
wire \mifu/_193_ ;
wire \mifu/_194_ ;
wire \mifu/_195_ ;
wire \mifu/_196_ ;
wire \mifu/_197_ ;
wire \mifu/_198_ ;
wire \mifu/_199_ ;
wire \mifu/_200_ ;
wire \mifu/_201_ ;
wire \mifu/_202_ ;
wire \mifu/_203_ ;
wire \mifu/_204_ ;
wire \mifu/_205_ ;
wire \mifu/_206_ ;
wire \mifu/_207_ ;
wire \mifu/_208_ ;
wire \mifu/_209_ ;
wire \mifu/_210_ ;
wire \mifu/_211_ ;
wire \mifu/_212_ ;
wire \mifu/_213_ ;
wire \mifu/_214_ ;
wire \mifu/_215_ ;
wire \mifu/_216_ ;
wire \mifu/_217_ ;
wire \mifu/_218_ ;
wire \mifu/_219_ ;
wire \mifu/_220_ ;
wire \mifu/_221_ ;
wire \mifu/_222_ ;
wire \mifu/_223_ ;
wire \mifu/wait_ready ;
wire \mlsu/_000_ ;
wire \mlsu/_001_ ;
wire \mlsu/_002_ ;
wire \mlsu/_003_ ;
wire \mlsu/_004_ ;
wire \mlsu/_005_ ;
wire \mlsu/_006_ ;
wire \mlsu/_007_ ;
wire \mlsu/_008_ ;
wire \mlsu/_009_ ;
wire \mlsu/_010_ ;
wire \mlsu/_011_ ;
wire \mlsu/_012_ ;
wire \mlsu/_013_ ;
wire \mlsu/_014_ ;
wire \mlsu/_015_ ;
wire \mlsu/_016_ ;
wire \mlsu/_017_ ;
wire \mlsu/_018_ ;
wire \mlsu/_019_ ;
wire \mlsu/_020_ ;
wire \mlsu/_021_ ;
wire \mlsu/_022_ ;
wire \mlsu/_023_ ;
wire \mlsu/_024_ ;
wire \mlsu/_025_ ;
wire \mlsu/_026_ ;
wire \mlsu/_027_ ;
wire \mlsu/_028_ ;
wire \mlsu/_029_ ;
wire \mlsu/_030_ ;
wire \mlsu/_031_ ;
wire \mlsu/_032_ ;
wire \mlsu/_033_ ;
wire \mlsu/_034_ ;
wire \mlsu/_035_ ;
wire \mlsu/_036_ ;
wire \mlsu/_037_ ;
wire \mlsu/_038_ ;
wire \mlsu/_039_ ;
wire \mlsu/_040_ ;
wire \mlsu/_041_ ;
wire \mlsu/_042_ ;
wire \mlsu/_043_ ;
wire \mlsu/_044_ ;
wire \mlsu/_045_ ;
wire \mlsu/_046_ ;
wire \mlsu/_047_ ;
wire \mlsu/_048_ ;
wire \mlsu/_049_ ;
wire \mlsu/_050_ ;
wire \mlsu/_051_ ;
wire \mlsu/_052_ ;
wire \mlsu/_053_ ;
wire \mlsu/_054_ ;
wire \mlsu/_055_ ;
wire \mlsu/_056_ ;
wire \mlsu/_057_ ;
wire \mlsu/_058_ ;
wire \mlsu/_059_ ;
wire \mlsu/_060_ ;
wire \mlsu/_061_ ;
wire \mlsu/_062_ ;
wire \mlsu/_063_ ;
wire \mlsu/_064_ ;
wire \mlsu/_065_ ;
wire \mlsu/_066_ ;
wire \mlsu/_067_ ;
wire \mlsu/_068_ ;
wire \mlsu/_069_ ;
wire \mlsu/_070_ ;
wire \mlsu/_071_ ;
wire \mlsu/_072_ ;
wire \mlsu/_073_ ;
wire \mlsu/_074_ ;
wire \mlsu/_075_ ;
wire \mlsu/_076_ ;
wire \mlsu/_077_ ;
wire \mlsu/_078_ ;
wire \mlsu/_079_ ;
wire \mlsu/_080_ ;
wire \mlsu/_081_ ;
wire \mlsu/_082_ ;
wire \mlsu/_083_ ;
wire \mlsu/_084_ ;
wire \mlsu/_085_ ;
wire \mlsu/_086_ ;
wire \mlsu/_087_ ;
wire \mlsu/_088_ ;
wire \mlsu/_089_ ;
wire \mlsu/_090_ ;
wire \mlsu/_091_ ;
wire \mlsu/_092_ ;
wire \mlsu/_093_ ;
wire \mlsu/_094_ ;
wire \mlsu/_095_ ;
wire \mlsu/_096_ ;
wire \mlsu/_097_ ;
wire \mlsu/_098_ ;
wire \mlsu/_099_ ;
wire \mlsu/_100_ ;
wire \mlsu/_101_ ;
wire \mlsu/_102_ ;
wire \mlsu/_103_ ;
wire \mlsu/_104_ ;
wire \mlsu/_105_ ;
wire \mlsu/_106_ ;
wire \mlsu/_107_ ;
wire \mlsu/_108_ ;
wire \mlsu/_109_ ;
wire \mlsu/_110_ ;
wire \mlsu/_111_ ;
wire \mlsu/_112_ ;
wire \mlsu/_113_ ;
wire \mlsu/_114_ ;
wire \mlsu/_115_ ;
wire \mlsu/_116_ ;
wire \mlsu/_117_ ;
wire \mlsu/_118_ ;
wire \mlsu/_119_ ;
wire \mlsu/_120_ ;
wire \mlsu/_121_ ;
wire \mlsu/_122_ ;
wire \mlsu/_123_ ;
wire \mlsu/_124_ ;
wire \mlsu/_125_ ;
wire \mlsu/_126_ ;
wire \mlsu/_127_ ;
wire \mlsu/_128_ ;
wire \mlsu/_129_ ;
wire \mlsu/_130_ ;
wire \mlsu/_131_ ;
wire \mlsu/_132_ ;
wire \mlsu/_133_ ;
wire \mlsu/_134_ ;
wire \mlsu/_135_ ;
wire \mlsu/_136_ ;
wire \mlsu/_137_ ;
wire \mlsu/_138_ ;
wire \mlsu/_139_ ;
wire \mlsu/_140_ ;
wire \mlsu/_141_ ;
wire \mlsu/_142_ ;
wire \mlsu/_143_ ;
wire \mlsu/_144_ ;
wire \mlsu/_145_ ;
wire \mlsu/_146_ ;
wire \mlsu/_147_ ;
wire \mlsu/_148_ ;
wire \mlsu/_149_ ;
wire \mlsu/_150_ ;
wire \mlsu/_151_ ;
wire \mlsu/_152_ ;
wire \mlsu/_153_ ;
wire \mlsu/_154_ ;
wire \mlsu/_155_ ;
wire \mlsu/_156_ ;
wire \mlsu/_157_ ;
wire \mlsu/_158_ ;
wire \mlsu/_159_ ;
wire \mlsu/_160_ ;
wire \mlsu/_161_ ;
wire \mlsu/_162_ ;
wire \mlsu/_163_ ;
wire \mlsu/_164_ ;
wire \mlsu/_165_ ;
wire \mlsu/_166_ ;
wire \mlsu/_167_ ;
wire \mlsu/_168_ ;
wire \mlsu/_169_ ;
wire \mlsu/_170_ ;
wire \mlsu/_171_ ;
wire \mlsu/_172_ ;
wire \mlsu/_173_ ;
wire \mlsu/_174_ ;
wire \mlsu/_175_ ;
wire \mlsu/_176_ ;
wire \mlsu/_177_ ;
wire \mlsu/_178_ ;
wire \mlsu/_179_ ;
wire \mlsu/_180_ ;
wire \mlsu/_181_ ;
wire \mlsu/_182_ ;
wire \mlsu/_183_ ;
wire \mlsu/_184_ ;
wire \mlsu/_185_ ;
wire \mlsu/_186_ ;
wire \mlsu/_187_ ;
wire \mlsu/_188_ ;
wire \mlsu/_189_ ;
wire \mlsu/_190_ ;
wire \mlsu/_191_ ;
wire \mlsu/_192_ ;
wire \mlsu/_193_ ;
wire \mlsu/_194_ ;
wire \mlsu/_195_ ;
wire \mlsu/_196_ ;
wire \mlsu/_197_ ;
wire \mlsu/_198_ ;
wire \mlsu/_199_ ;
wire \mlsu/_200_ ;
wire \mlsu/_201_ ;
wire \mlsu/_202_ ;
wire \mlsu/_203_ ;
wire \mlsu/_204_ ;
wire \mlsu/_205_ ;
wire \mlsu/_206_ ;
wire \mlsu/_207_ ;
wire \mlsu/_208_ ;
wire \mlsu/_209_ ;
wire \mlsu/_210_ ;
wire \mlsu/_211_ ;
wire \mlsu/_212_ ;
wire \mlsu/_213_ ;
wire \mlsu/_214_ ;
wire \mlsu/_215_ ;
wire \mlsu/_216_ ;
wire \mlsu/_217_ ;
wire \mlsu/_218_ ;
wire \mlsu/_219_ ;
wire \mlsu/_220_ ;
wire \mlsu/_221_ ;
wire \mlsu/_222_ ;
wire \mlsu/_223_ ;
wire \mlsu/_224_ ;
wire \mlsu/_225_ ;
wire \mlsu/_226_ ;
wire \mlsu/_227_ ;
wire \mlsu/_228_ ;
wire \mlsu/_229_ ;
wire \mlsu/_230_ ;
wire \mlsu/_231_ ;
wire \mlsu/_232_ ;
wire \mlsu/_233_ ;
wire \mlsu/_234_ ;
wire \mlsu/_235_ ;
wire \mlsu/_236_ ;
wire \mlsu/_237_ ;
wire \mlsu/_238_ ;
wire \mlsu/_239_ ;
wire \mlsu/_240_ ;
wire \mlsu/_241_ ;
wire \mlsu/_242_ ;
wire \mlsu/_243_ ;
wire \mlsu/_244_ ;
wire \mlsu/_245_ ;
wire \mlsu/_246_ ;
wire \mlsu/_247_ ;
wire \mlsu/_248_ ;
wire \mlsu/_249_ ;
wire \mlsu/_250_ ;
wire \mlsu/_251_ ;
wire \mlsu/_252_ ;
wire \mlsu/_253_ ;
wire \mlsu/_254_ ;
wire \mlsu/_255_ ;
wire \mlsu/_256_ ;
wire \mlsu/_257_ ;
wire \mlsu/_258_ ;
wire \mlsu/_259_ ;
wire \mlsu/_260_ ;
wire \mlsu/_261_ ;
wire \mlsu/_262_ ;
wire \mlsu/_263_ ;
wire \mlsu/_264_ ;
wire \mlsu/_265_ ;
wire \mlsu/_266_ ;
wire \mlsu/_267_ ;
wire \mlsu/_268_ ;
wire \mlsu/_269_ ;
wire \mlsu/_rdata[0] ;
wire \mlsu/_rdata[10] ;
wire \mlsu/_rdata[11] ;
wire \mlsu/_rdata[12] ;
wire \mlsu/_rdata[13] ;
wire \mlsu/_rdata[14] ;
wire \mlsu/_rdata[15] ;
wire \mlsu/_rdata[16] ;
wire \mlsu/_rdata[17] ;
wire \mlsu/_rdata[18] ;
wire \mlsu/_rdata[19] ;
wire \mlsu/_rdata[1] ;
wire \mlsu/_rdata[20] ;
wire \mlsu/_rdata[21] ;
wire \mlsu/_rdata[22] ;
wire \mlsu/_rdata[23] ;
wire \mlsu/_rdata[24] ;
wire \mlsu/_rdata[25] ;
wire \mlsu/_rdata[26] ;
wire \mlsu/_rdata[27] ;
wire \mlsu/_rdata[28] ;
wire \mlsu/_rdata[29] ;
wire \mlsu/_rdata[2] ;
wire \mlsu/_rdata[30] ;
wire \mlsu/_rdata[31] ;
wire \mlsu/_rdata[3] ;
wire \mlsu/_rdata[4] ;
wire \mlsu/_rdata[5] ;
wire \mlsu/_rdata[6] ;
wire \mlsu/_rdata[7] ;
wire \mlsu/_rdata[8] ;
wire \mlsu/_rdata[9] ;
wire \mlsu/write_wait_ready ;
wire \mpc/_000_ ;
wire \mpc/_001_ ;
wire \mpc/_002_ ;
wire \mpc/_003_ ;
wire \mpc/_004_ ;
wire \mpc/_005_ ;
wire \mpc/_006_ ;
wire \mpc/_007_ ;
wire \mpc/_008_ ;
wire \mpc/_009_ ;
wire \mpc/_010_ ;
wire \mpc/_011_ ;
wire \mpc/_012_ ;
wire \mpc/_013_ ;
wire \mpc/_014_ ;
wire \mpc/_015_ ;
wire \mpc/_016_ ;
wire \mpc/_017_ ;
wire \mpc/_018_ ;
wire \mpc/_019_ ;
wire \mpc/_020_ ;
wire \mpc/_021_ ;
wire \mpc/_022_ ;
wire \mpc/_023_ ;
wire \mpc/_024_ ;
wire \mpc/_025_ ;
wire \mpc/_026_ ;
wire \mpc/_027_ ;
wire \mpc/_028_ ;
wire \mpc/_029_ ;
wire \mpc/_030_ ;
wire \mpc/_031_ ;
wire \mpc/_032_ ;
wire \mpc/_033_ ;
wire \mpc/_034_ ;
wire \mpc/_035_ ;
wire \mpc/_036_ ;
wire \mpc/_037_ ;
wire \mpc/_038_ ;
wire \mpc/_039_ ;
wire \mpc/_040_ ;
wire \mpc/_041_ ;
wire \mpc/_042_ ;
wire \mpc/_043_ ;
wire \mpc/_044_ ;
wire \mpc/_045_ ;
wire \mpc/_046_ ;
wire \mpc/_047_ ;
wire \mpc/_048_ ;
wire \mpc/_049_ ;
wire \mpc/_050_ ;
wire \mpc/_051_ ;
wire \mpc/_052_ ;
wire \mpc/_053_ ;
wire \mpc/_054_ ;
wire \mpc/_055_ ;
wire \mpc/_056_ ;
wire \mpc/_057_ ;
wire \mpc/_058_ ;
wire \mpc/_059_ ;
wire \mpc/_060_ ;
wire \mpc/_061_ ;
wire \mpc/_062_ ;
wire \mpc/_063_ ;
wire \mpc/_064_ ;
wire \mpc/_065_ ;
wire \mpc/_066_ ;
wire \mpc/_067_ ;
wire \mpc/_068_ ;
wire \mpc/_069_ ;
wire \mpc/_070_ ;
wire \mpc/_071_ ;
wire \mpc/_072_ ;
wire \mpc/_073_ ;
wire \mpc/_074_ ;
wire \mpc/_075_ ;
wire \mpc/_076_ ;
wire \mpc/_077_ ;
wire \mpc/_078_ ;
wire \mpc/_079_ ;
wire \mpc/_080_ ;
wire \mpc/_081_ ;
wire \mpc/_082_ ;
wire \mpc/_083_ ;
wire \mpc/_084_ ;
wire \mpc/_085_ ;
wire \mpc/_086_ ;
wire \mpc/_087_ ;
wire \mpc/_088_ ;
wire \mpc/_089_ ;
wire \mpc/_090_ ;
wire \mpc/_091_ ;
wire \mpc/_092_ ;
wire \mpc/_093_ ;
wire \mpc/_094_ ;
wire \mpc/_095_ ;
wire \mpc/_096_ ;
wire \mpc/_097_ ;
wire \mpc/_098_ ;
wire \mpc/_099_ ;
wire \mpc/_100_ ;
wire \mpc/_101_ ;
wire \mpc/_102_ ;
wire \mpc/_103_ ;
wire \mpc/_104_ ;
wire \mpc/_105_ ;
wire \mpc/_106_ ;
wire \mpc/_107_ ;
wire \mpc/_108_ ;
wire \mpc/_109_ ;
wire \mpc/_110_ ;
wire \mpc/_111_ ;
wire \mpc/_112_ ;
wire \mpc/_113_ ;
wire \mpc/_114_ ;
wire \mpc/_115_ ;
wire \mpc/_116_ ;
wire \mpc/_117_ ;
wire \mpc/_118_ ;
wire \mpc/_119_ ;
wire \mpc/_120_ ;
wire \mpc/_121_ ;
wire \mpc/_122_ ;
wire \mpc/_123_ ;
wire \mpc/_124_ ;
wire \mpc/_125_ ;
wire \mpc/_126_ ;
wire \mpc/_127_ ;
wire \mpc/_128_ ;
wire \mpc/_129_ ;
wire \mpc/_130_ ;
wire \mpc/_131_ ;
wire \mpc/_132_ ;
wire \mpc/_133_ ;
wire \mpc/_134_ ;
wire \mpc/_135_ ;
wire \mpc/_136_ ;
wire \mpc/_137_ ;
wire \mpc/_138_ ;
wire \mpc/_139_ ;
wire \mpc/_140_ ;
wire \mpc/_141_ ;
wire \mpc/_142_ ;
wire \mpc/_143_ ;
wire \mpc/_144_ ;
wire \mpc/_145_ ;
wire \mpc/_146_ ;
wire \mpc/_147_ ;
wire \mpc/_148_ ;
wire \mpc/_149_ ;
wire \mpc/_150_ ;
wire \mpc/_151_ ;
wire \mpc/_152_ ;
wire \mpc/_153_ ;
wire \mpc/_154_ ;
wire \mpc/_155_ ;
wire \mpc/_156_ ;
wire \mpc/_157_ ;
wire \mpc/_158_ ;
wire \mpc/_159_ ;
wire \mpc/_160_ ;
wire \mpc/_161_ ;
wire \mpc/_162_ ;
wire \mpc/_163_ ;
wire \mpc/_164_ ;
wire \mpc/_165_ ;
wire \mpc/_166_ ;
wire \mpc/_167_ ;
wire \mpc/_168_ ;
wire \mpc/_169_ ;
wire \mpc/_170_ ;
wire \mpc/_171_ ;
wire \mpc/_172_ ;
wire \mpc/_173_ ;
wire \mpc/_174_ ;
wire \mpc/_175_ ;
wire \mpc/_176_ ;
wire \mpc/_177_ ;
wire \mpc/_178_ ;
wire \mpc/_179_ ;
wire \mpc/_180_ ;
wire \mpc/_181_ ;
wire \mpc/_182_ ;
wire \mpc/_183_ ;
wire \mpc/_184_ ;
wire \mpc/_185_ ;
wire \mpc/_186_ ;
wire \mpc/_187_ ;
wire \mpc/_188_ ;
wire \mpc/_189_ ;
wire \mpc/_190_ ;
wire \mpc/_191_ ;
wire \mpc/_192_ ;
wire \mpc/_193_ ;
wire \mpc/_194_ ;
wire \mpc/_195_ ;
wire \mpc/_196_ ;
wire \mpc/_197_ ;
wire \mpc/_198_ ;
wire \mpc/_199_ ;
wire \mpc/_200_ ;
wire \mpc/_201_ ;
wire \mpc/_202_ ;
wire \mpc/_203_ ;
wire \mpc/_204_ ;
wire \mpc/_205_ ;
wire \mpc/_206_ ;
wire \mpc/_207_ ;
wire \mpc/_208_ ;
wire \mpc/_209_ ;
wire \mpc/_210_ ;
wire \mpc/_211_ ;
wire \mpc/_212_ ;
wire \mpc/_213_ ;
wire \mpc/_214_ ;
wire \mpc/_215_ ;
wire \mpc/_216_ ;
wire \mpc/_217_ ;
wire \mpc/_218_ ;
wire \mpc/_219_ ;
wire \mpc/_220_ ;
wire \mpc/_221_ ;
wire \mpc/_222_ ;
wire \mpc/_223_ ;
wire \mpc/_224_ ;
wire \mpc/_225_ ;
wire \mpc/_226_ ;
wire \mpc/_227_ ;
wire \mpc/_228_ ;
wire \mpc/_229_ ;
wire \mpc/_230_ ;
wire \mpc/_231_ ;
wire \mpc/_232_ ;
wire \mpc/_233_ ;
wire \mpc/_234_ ;
wire \mpc/_235_ ;
wire \mpc/_236_ ;
wire \mpc/_237_ ;
wire \mpc/_238_ ;
wire \mpc/_239_ ;
wire \mpc/_240_ ;
wire \mpc/_241_ ;
wire \mpc/_242_ ;
wire \mpc/_243_ ;
wire \mpc/_244_ ;
wire \mpc/_245_ ;
wire \mpc/_246_ ;
wire \mpc/_247_ ;
wire \mpc/_248_ ;
wire \mpc/_249_ ;
wire \mpc/_250_ ;
wire \mpc/_251_ ;
wire \mpc/_252_ ;
wire \mpc/_253_ ;
wire \mpc/_254_ ;
wire \mpc/_255_ ;
wire \mpc/_256_ ;
wire \mpc/_257_ ;
wire \mpc/_258_ ;
wire \mpc/_259_ ;
wire \mpc/_260_ ;
wire \mpc/_261_ ;
wire \mpc/_262_ ;
wire \mpc/_263_ ;
wire \mpc/_264_ ;
wire \mpc/_265_ ;
wire \mpc/_266_ ;
wire \mpc/_267_ ;
wire \mpc/_268_ ;
wire \mpc/_269_ ;
wire \mpc/_270_ ;
wire \mpc/_271_ ;
wire \mpc/_272_ ;
wire \mpc/_273_ ;
wire \mpc/_274_ ;
wire \mpc/_275_ ;
wire \mpc/_276_ ;
wire \mpc/_277_ ;
wire \mpc/_278_ ;
wire \mpc/_279_ ;
wire \mpc/_280_ ;
wire \mpc/_281_ ;
wire \mpc/_282_ ;
wire \mpc/_283_ ;
wire \mpc/_284_ ;
wire \mpc/_285_ ;
wire \mpc/_286_ ;
wire \mpc/_287_ ;
wire \mpc/_288_ ;
wire \mpc/_289_ ;
wire \mpc/_290_ ;
wire \mpc/_291_ ;
wire \mpc/_292_ ;
wire \mpc/_293_ ;
wire \mpc/_294_ ;
wire \mpc/_295_ ;
wire \mpc/_296_ ;
wire \mpc/_297_ ;
wire \mpc/_298_ ;
wire \mpc/_299_ ;
wire \mpc/_300_ ;
wire \mpc/_301_ ;
wire \mpc/_302_ ;
wire \mpc/_303_ ;
wire \mpc/_304_ ;
wire \mpc/_305_ ;
wire \mpc/_306_ ;
wire \mpc/_307_ ;
wire \mpc/_308_ ;
wire \mpc/_309_ ;
wire \mpc/_310_ ;
wire \mpc/_311_ ;
wire \mpc/_312_ ;
wire \mpc/_313_ ;
wire \mpc/_314_ ;
wire \mpc/_315_ ;
wire \mpc/_316_ ;
wire \mpc/_317_ ;
wire \mpc/_318_ ;
wire \mpc/_319_ ;
wire \mpc/_320_ ;
wire \mpc/_321_ ;
wire \mpc/_322_ ;
wire \mpc/_323_ ;
wire \mpc/_324_ ;
wire \mpc/_325_ ;
wire \mpc/_326_ ;
wire \mreg/_00000_ ;
wire \mreg/_00001_ ;
wire \mreg/_00002_ ;
wire \mreg/_00003_ ;
wire \mreg/_00004_ ;
wire \mreg/_00005_ ;
wire \mreg/_00006_ ;
wire \mreg/_00007_ ;
wire \mreg/_00008_ ;
wire \mreg/_00009_ ;
wire \mreg/_00010_ ;
wire \mreg/_00011_ ;
wire \mreg/_00012_ ;
wire \mreg/_00013_ ;
wire \mreg/_00014_ ;
wire \mreg/_00015_ ;
wire \mreg/_00016_ ;
wire \mreg/_00017_ ;
wire \mreg/_00018_ ;
wire \mreg/_00019_ ;
wire \mreg/_00020_ ;
wire \mreg/_00021_ ;
wire \mreg/_00022_ ;
wire \mreg/_00023_ ;
wire \mreg/_00024_ ;
wire \mreg/_00025_ ;
wire \mreg/_00026_ ;
wire \mreg/_00027_ ;
wire \mreg/_00028_ ;
wire \mreg/_00029_ ;
wire \mreg/_00030_ ;
wire \mreg/_00031_ ;
wire \mreg/_00032_ ;
wire \mreg/_00033_ ;
wire \mreg/_00034_ ;
wire \mreg/_00035_ ;
wire \mreg/_00036_ ;
wire \mreg/_00037_ ;
wire \mreg/_00038_ ;
wire \mreg/_00039_ ;
wire \mreg/_00040_ ;
wire \mreg/_00041_ ;
wire \mreg/_00042_ ;
wire \mreg/_00043_ ;
wire \mreg/_00044_ ;
wire \mreg/_00045_ ;
wire \mreg/_00046_ ;
wire \mreg/_00047_ ;
wire \mreg/_00048_ ;
wire \mreg/_00049_ ;
wire \mreg/_00050_ ;
wire \mreg/_00051_ ;
wire \mreg/_00052_ ;
wire \mreg/_00053_ ;
wire \mreg/_00054_ ;
wire \mreg/_00055_ ;
wire \mreg/_00056_ ;
wire \mreg/_00057_ ;
wire \mreg/_00058_ ;
wire \mreg/_00059_ ;
wire \mreg/_00060_ ;
wire \mreg/_00061_ ;
wire \mreg/_00062_ ;
wire \mreg/_00063_ ;
wire \mreg/_00064_ ;
wire \mreg/_00065_ ;
wire \mreg/_00066_ ;
wire \mreg/_00067_ ;
wire \mreg/_00068_ ;
wire \mreg/_00069_ ;
wire \mreg/_00070_ ;
wire \mreg/_00071_ ;
wire \mreg/_00072_ ;
wire \mreg/_00073_ ;
wire \mreg/_00074_ ;
wire \mreg/_00075_ ;
wire \mreg/_00076_ ;
wire \mreg/_00077_ ;
wire \mreg/_00078_ ;
wire \mreg/_00079_ ;
wire \mreg/_00080_ ;
wire \mreg/_00081_ ;
wire \mreg/_00082_ ;
wire \mreg/_00083_ ;
wire \mreg/_00084_ ;
wire \mreg/_00085_ ;
wire \mreg/_00086_ ;
wire \mreg/_00087_ ;
wire \mreg/_00088_ ;
wire \mreg/_00089_ ;
wire \mreg/_00090_ ;
wire \mreg/_00091_ ;
wire \mreg/_00092_ ;
wire \mreg/_00093_ ;
wire \mreg/_00094_ ;
wire \mreg/_00095_ ;
wire \mreg/_00096_ ;
wire \mreg/_00097_ ;
wire \mreg/_00098_ ;
wire \mreg/_00099_ ;
wire \mreg/_00100_ ;
wire \mreg/_00101_ ;
wire \mreg/_00102_ ;
wire \mreg/_00103_ ;
wire \mreg/_00104_ ;
wire \mreg/_00105_ ;
wire \mreg/_00106_ ;
wire \mreg/_00107_ ;
wire \mreg/_00108_ ;
wire \mreg/_00109_ ;
wire \mreg/_00110_ ;
wire \mreg/_00111_ ;
wire \mreg/_00112_ ;
wire \mreg/_00113_ ;
wire \mreg/_00114_ ;
wire \mreg/_00115_ ;
wire \mreg/_00116_ ;
wire \mreg/_00117_ ;
wire \mreg/_00118_ ;
wire \mreg/_00119_ ;
wire \mreg/_00120_ ;
wire \mreg/_00121_ ;
wire \mreg/_00122_ ;
wire \mreg/_00123_ ;
wire \mreg/_00124_ ;
wire \mreg/_00125_ ;
wire \mreg/_00126_ ;
wire \mreg/_00127_ ;
wire \mreg/_00128_ ;
wire \mreg/_00129_ ;
wire \mreg/_00130_ ;
wire \mreg/_00131_ ;
wire \mreg/_00132_ ;
wire \mreg/_00133_ ;
wire \mreg/_00134_ ;
wire \mreg/_00135_ ;
wire \mreg/_00136_ ;
wire \mreg/_00137_ ;
wire \mreg/_00138_ ;
wire \mreg/_00139_ ;
wire \mreg/_00140_ ;
wire \mreg/_00141_ ;
wire \mreg/_00142_ ;
wire \mreg/_00143_ ;
wire \mreg/_00144_ ;
wire \mreg/_00145_ ;
wire \mreg/_00146_ ;
wire \mreg/_00147_ ;
wire \mreg/_00148_ ;
wire \mreg/_00149_ ;
wire \mreg/_00150_ ;
wire \mreg/_00151_ ;
wire \mreg/_00152_ ;
wire \mreg/_00153_ ;
wire \mreg/_00154_ ;
wire \mreg/_00155_ ;
wire \mreg/_00156_ ;
wire \mreg/_00157_ ;
wire \mreg/_00158_ ;
wire \mreg/_00159_ ;
wire \mreg/_00160_ ;
wire \mreg/_00161_ ;
wire \mreg/_00162_ ;
wire \mreg/_00163_ ;
wire \mreg/_00164_ ;
wire \mreg/_00165_ ;
wire \mreg/_00166_ ;
wire \mreg/_00167_ ;
wire \mreg/_00168_ ;
wire \mreg/_00169_ ;
wire \mreg/_00170_ ;
wire \mreg/_00171_ ;
wire \mreg/_00172_ ;
wire \mreg/_00173_ ;
wire \mreg/_00174_ ;
wire \mreg/_00175_ ;
wire \mreg/_00176_ ;
wire \mreg/_00177_ ;
wire \mreg/_00178_ ;
wire \mreg/_00179_ ;
wire \mreg/_00180_ ;
wire \mreg/_00181_ ;
wire \mreg/_00182_ ;
wire \mreg/_00183_ ;
wire \mreg/_00184_ ;
wire \mreg/_00185_ ;
wire \mreg/_00186_ ;
wire \mreg/_00187_ ;
wire \mreg/_00188_ ;
wire \mreg/_00189_ ;
wire \mreg/_00190_ ;
wire \mreg/_00191_ ;
wire \mreg/_00192_ ;
wire \mreg/_00193_ ;
wire \mreg/_00194_ ;
wire \mreg/_00195_ ;
wire \mreg/_00196_ ;
wire \mreg/_00197_ ;
wire \mreg/_00198_ ;
wire \mreg/_00199_ ;
wire \mreg/_00200_ ;
wire \mreg/_00201_ ;
wire \mreg/_00202_ ;
wire \mreg/_00203_ ;
wire \mreg/_00204_ ;
wire \mreg/_00205_ ;
wire \mreg/_00206_ ;
wire \mreg/_00207_ ;
wire \mreg/_00208_ ;
wire \mreg/_00209_ ;
wire \mreg/_00210_ ;
wire \mreg/_00211_ ;
wire \mreg/_00212_ ;
wire \mreg/_00213_ ;
wire \mreg/_00214_ ;
wire \mreg/_00215_ ;
wire \mreg/_00216_ ;
wire \mreg/_00217_ ;
wire \mreg/_00218_ ;
wire \mreg/_00219_ ;
wire \mreg/_00220_ ;
wire \mreg/_00221_ ;
wire \mreg/_00222_ ;
wire \mreg/_00223_ ;
wire \mreg/_00224_ ;
wire \mreg/_00225_ ;
wire \mreg/_00226_ ;
wire \mreg/_00227_ ;
wire \mreg/_00228_ ;
wire \mreg/_00229_ ;
wire \mreg/_00230_ ;
wire \mreg/_00231_ ;
wire \mreg/_00232_ ;
wire \mreg/_00233_ ;
wire \mreg/_00234_ ;
wire \mreg/_00235_ ;
wire \mreg/_00236_ ;
wire \mreg/_00237_ ;
wire \mreg/_00238_ ;
wire \mreg/_00239_ ;
wire \mreg/_00240_ ;
wire \mreg/_00241_ ;
wire \mreg/_00242_ ;
wire \mreg/_00243_ ;
wire \mreg/_00244_ ;
wire \mreg/_00245_ ;
wire \mreg/_00246_ ;
wire \mreg/_00247_ ;
wire \mreg/_00248_ ;
wire \mreg/_00249_ ;
wire \mreg/_00250_ ;
wire \mreg/_00251_ ;
wire \mreg/_00252_ ;
wire \mreg/_00253_ ;
wire \mreg/_00254_ ;
wire \mreg/_00255_ ;
wire \mreg/_00256_ ;
wire \mreg/_00257_ ;
wire \mreg/_00258_ ;
wire \mreg/_00259_ ;
wire \mreg/_00260_ ;
wire \mreg/_00261_ ;
wire \mreg/_00262_ ;
wire \mreg/_00263_ ;
wire \mreg/_00264_ ;
wire \mreg/_00265_ ;
wire \mreg/_00266_ ;
wire \mreg/_00267_ ;
wire \mreg/_00268_ ;
wire \mreg/_00269_ ;
wire \mreg/_00270_ ;
wire \mreg/_00271_ ;
wire \mreg/_00272_ ;
wire \mreg/_00273_ ;
wire \mreg/_00274_ ;
wire \mreg/_00275_ ;
wire \mreg/_00276_ ;
wire \mreg/_00277_ ;
wire \mreg/_00278_ ;
wire \mreg/_00279_ ;
wire \mreg/_00280_ ;
wire \mreg/_00281_ ;
wire \mreg/_00282_ ;
wire \mreg/_00283_ ;
wire \mreg/_00284_ ;
wire \mreg/_00285_ ;
wire \mreg/_00286_ ;
wire \mreg/_00287_ ;
wire \mreg/_00288_ ;
wire \mreg/_00289_ ;
wire \mreg/_00290_ ;
wire \mreg/_00291_ ;
wire \mreg/_00292_ ;
wire \mreg/_00293_ ;
wire \mreg/_00294_ ;
wire \mreg/_00295_ ;
wire \mreg/_00296_ ;
wire \mreg/_00297_ ;
wire \mreg/_00298_ ;
wire \mreg/_00299_ ;
wire \mreg/_00300_ ;
wire \mreg/_00301_ ;
wire \mreg/_00302_ ;
wire \mreg/_00303_ ;
wire \mreg/_00304_ ;
wire \mreg/_00305_ ;
wire \mreg/_00306_ ;
wire \mreg/_00307_ ;
wire \mreg/_00308_ ;
wire \mreg/_00309_ ;
wire \mreg/_00310_ ;
wire \mreg/_00311_ ;
wire \mreg/_00312_ ;
wire \mreg/_00313_ ;
wire \mreg/_00314_ ;
wire \mreg/_00315_ ;
wire \mreg/_00316_ ;
wire \mreg/_00317_ ;
wire \mreg/_00318_ ;
wire \mreg/_00319_ ;
wire \mreg/_00320_ ;
wire \mreg/_00321_ ;
wire \mreg/_00322_ ;
wire \mreg/_00323_ ;
wire \mreg/_00324_ ;
wire \mreg/_00325_ ;
wire \mreg/_00326_ ;
wire \mreg/_00327_ ;
wire \mreg/_00328_ ;
wire \mreg/_00329_ ;
wire \mreg/_00330_ ;
wire \mreg/_00331_ ;
wire \mreg/_00332_ ;
wire \mreg/_00333_ ;
wire \mreg/_00334_ ;
wire \mreg/_00335_ ;
wire \mreg/_00336_ ;
wire \mreg/_00337_ ;
wire \mreg/_00338_ ;
wire \mreg/_00339_ ;
wire \mreg/_00340_ ;
wire \mreg/_00341_ ;
wire \mreg/_00342_ ;
wire \mreg/_00343_ ;
wire \mreg/_00344_ ;
wire \mreg/_00345_ ;
wire \mreg/_00346_ ;
wire \mreg/_00347_ ;
wire \mreg/_00348_ ;
wire \mreg/_00349_ ;
wire \mreg/_00350_ ;
wire \mreg/_00351_ ;
wire \mreg/_00352_ ;
wire \mreg/_00353_ ;
wire \mreg/_00354_ ;
wire \mreg/_00355_ ;
wire \mreg/_00356_ ;
wire \mreg/_00357_ ;
wire \mreg/_00358_ ;
wire \mreg/_00359_ ;
wire \mreg/_00360_ ;
wire \mreg/_00361_ ;
wire \mreg/_00362_ ;
wire \mreg/_00363_ ;
wire \mreg/_00364_ ;
wire \mreg/_00365_ ;
wire \mreg/_00366_ ;
wire \mreg/_00367_ ;
wire \mreg/_00368_ ;
wire \mreg/_00369_ ;
wire \mreg/_00370_ ;
wire \mreg/_00371_ ;
wire \mreg/_00372_ ;
wire \mreg/_00373_ ;
wire \mreg/_00374_ ;
wire \mreg/_00375_ ;
wire \mreg/_00376_ ;
wire \mreg/_00377_ ;
wire \mreg/_00378_ ;
wire \mreg/_00379_ ;
wire \mreg/_00380_ ;
wire \mreg/_00381_ ;
wire \mreg/_00382_ ;
wire \mreg/_00383_ ;
wire \mreg/_00384_ ;
wire \mreg/_00385_ ;
wire \mreg/_00386_ ;
wire \mreg/_00387_ ;
wire \mreg/_00388_ ;
wire \mreg/_00389_ ;
wire \mreg/_00390_ ;
wire \mreg/_00391_ ;
wire \mreg/_00392_ ;
wire \mreg/_00393_ ;
wire \mreg/_00394_ ;
wire \mreg/_00395_ ;
wire \mreg/_00396_ ;
wire \mreg/_00397_ ;
wire \mreg/_00398_ ;
wire \mreg/_00399_ ;
wire \mreg/_00400_ ;
wire \mreg/_00401_ ;
wire \mreg/_00402_ ;
wire \mreg/_00403_ ;
wire \mreg/_00404_ ;
wire \mreg/_00405_ ;
wire \mreg/_00406_ ;
wire \mreg/_00407_ ;
wire \mreg/_00408_ ;
wire \mreg/_00409_ ;
wire \mreg/_00410_ ;
wire \mreg/_00411_ ;
wire \mreg/_00412_ ;
wire \mreg/_00413_ ;
wire \mreg/_00414_ ;
wire \mreg/_00415_ ;
wire \mreg/_00416_ ;
wire \mreg/_00417_ ;
wire \mreg/_00418_ ;
wire \mreg/_00419_ ;
wire \mreg/_00420_ ;
wire \mreg/_00421_ ;
wire \mreg/_00422_ ;
wire \mreg/_00423_ ;
wire \mreg/_00424_ ;
wire \mreg/_00425_ ;
wire \mreg/_00426_ ;
wire \mreg/_00427_ ;
wire \mreg/_00428_ ;
wire \mreg/_00429_ ;
wire \mreg/_00430_ ;
wire \mreg/_00431_ ;
wire \mreg/_00432_ ;
wire \mreg/_00433_ ;
wire \mreg/_00434_ ;
wire \mreg/_00435_ ;
wire \mreg/_00436_ ;
wire \mreg/_00437_ ;
wire \mreg/_00438_ ;
wire \mreg/_00439_ ;
wire \mreg/_00440_ ;
wire \mreg/_00441_ ;
wire \mreg/_00442_ ;
wire \mreg/_00443_ ;
wire \mreg/_00444_ ;
wire \mreg/_00445_ ;
wire \mreg/_00446_ ;
wire \mreg/_00447_ ;
wire \mreg/_00448_ ;
wire \mreg/_00449_ ;
wire \mreg/_00450_ ;
wire \mreg/_00451_ ;
wire \mreg/_00452_ ;
wire \mreg/_00453_ ;
wire \mreg/_00454_ ;
wire \mreg/_00455_ ;
wire \mreg/_00456_ ;
wire \mreg/_00457_ ;
wire \mreg/_00458_ ;
wire \mreg/_00459_ ;
wire \mreg/_00460_ ;
wire \mreg/_00461_ ;
wire \mreg/_00462_ ;
wire \mreg/_00463_ ;
wire \mreg/_00464_ ;
wire \mreg/_00465_ ;
wire \mreg/_00466_ ;
wire \mreg/_00467_ ;
wire \mreg/_00468_ ;
wire \mreg/_00469_ ;
wire \mreg/_00470_ ;
wire \mreg/_00471_ ;
wire \mreg/_00472_ ;
wire \mreg/_00473_ ;
wire \mreg/_00474_ ;
wire \mreg/_00475_ ;
wire \mreg/_00476_ ;
wire \mreg/_00477_ ;
wire \mreg/_00478_ ;
wire \mreg/_00479_ ;
wire \mreg/_00480_ ;
wire \mreg/_00481_ ;
wire \mreg/_00482_ ;
wire \mreg/_00483_ ;
wire \mreg/_00484_ ;
wire \mreg/_00485_ ;
wire \mreg/_00486_ ;
wire \mreg/_00487_ ;
wire \mreg/_00488_ ;
wire \mreg/_00489_ ;
wire \mreg/_00490_ ;
wire \mreg/_00491_ ;
wire \mreg/_00492_ ;
wire \mreg/_00493_ ;
wire \mreg/_00494_ ;
wire \mreg/_00495_ ;
wire \mreg/_00496_ ;
wire \mreg/_00497_ ;
wire \mreg/_00498_ ;
wire \mreg/_00499_ ;
wire \mreg/_00500_ ;
wire \mreg/_00501_ ;
wire \mreg/_00502_ ;
wire \mreg/_00503_ ;
wire \mreg/_00504_ ;
wire \mreg/_00505_ ;
wire \mreg/_00506_ ;
wire \mreg/_00507_ ;
wire \mreg/_00508_ ;
wire \mreg/_00509_ ;
wire \mreg/_00510_ ;
wire \mreg/_00511_ ;
wire \mreg/_00512_ ;
wire \mreg/_00513_ ;
wire \mreg/_00514_ ;
wire \mreg/_00515_ ;
wire \mreg/_00516_ ;
wire \mreg/_00517_ ;
wire \mreg/_00518_ ;
wire \mreg/_00519_ ;
wire \mreg/_00520_ ;
wire \mreg/_00521_ ;
wire \mreg/_00522_ ;
wire \mreg/_00523_ ;
wire \mreg/_00524_ ;
wire \mreg/_00525_ ;
wire \mreg/_00526_ ;
wire \mreg/_00527_ ;
wire \mreg/_00528_ ;
wire \mreg/_00529_ ;
wire \mreg/_00530_ ;
wire \mreg/_00531_ ;
wire \mreg/_00532_ ;
wire \mreg/_00533_ ;
wire \mreg/_00534_ ;
wire \mreg/_00535_ ;
wire \mreg/_00536_ ;
wire \mreg/_00537_ ;
wire \mreg/_00538_ ;
wire \mreg/_00539_ ;
wire \mreg/_00540_ ;
wire \mreg/_00541_ ;
wire \mreg/_00542_ ;
wire \mreg/_00543_ ;
wire \mreg/_00544_ ;
wire \mreg/_00545_ ;
wire \mreg/_00546_ ;
wire \mreg/_00547_ ;
wire \mreg/_00548_ ;
wire \mreg/_00549_ ;
wire \mreg/_00550_ ;
wire \mreg/_00551_ ;
wire \mreg/_00552_ ;
wire \mreg/_00553_ ;
wire \mreg/_00554_ ;
wire \mreg/_00555_ ;
wire \mreg/_00556_ ;
wire \mreg/_00557_ ;
wire \mreg/_00558_ ;
wire \mreg/_00559_ ;
wire \mreg/_00560_ ;
wire \mreg/_00561_ ;
wire \mreg/_00562_ ;
wire \mreg/_00563_ ;
wire \mreg/_00564_ ;
wire \mreg/_00565_ ;
wire \mreg/_00566_ ;
wire \mreg/_00567_ ;
wire \mreg/_00568_ ;
wire \mreg/_00569_ ;
wire \mreg/_00570_ ;
wire \mreg/_00571_ ;
wire \mreg/_00572_ ;
wire \mreg/_00573_ ;
wire \mreg/_00574_ ;
wire \mreg/_00575_ ;
wire \mreg/_00576_ ;
wire \mreg/_00577_ ;
wire \mreg/_00578_ ;
wire \mreg/_00579_ ;
wire \mreg/_00580_ ;
wire \mreg/_00581_ ;
wire \mreg/_00582_ ;
wire \mreg/_00583_ ;
wire \mreg/_00584_ ;
wire \mreg/_00585_ ;
wire \mreg/_00586_ ;
wire \mreg/_00587_ ;
wire \mreg/_00588_ ;
wire \mreg/_00589_ ;
wire \mreg/_00590_ ;
wire \mreg/_00591_ ;
wire \mreg/_00592_ ;
wire \mreg/_00593_ ;
wire \mreg/_00594_ ;
wire \mreg/_00595_ ;
wire \mreg/_00596_ ;
wire \mreg/_00597_ ;
wire \mreg/_00598_ ;
wire \mreg/_00599_ ;
wire \mreg/_00600_ ;
wire \mreg/_00601_ ;
wire \mreg/_00602_ ;
wire \mreg/_00603_ ;
wire \mreg/_00604_ ;
wire \mreg/_00605_ ;
wire \mreg/_00606_ ;
wire \mreg/_00607_ ;
wire \mreg/_00608_ ;
wire \mreg/_00609_ ;
wire \mreg/_00610_ ;
wire \mreg/_00611_ ;
wire \mreg/_00612_ ;
wire \mreg/_00613_ ;
wire \mreg/_00614_ ;
wire \mreg/_00615_ ;
wire \mreg/_00616_ ;
wire \mreg/_00617_ ;
wire \mreg/_00618_ ;
wire \mreg/_00619_ ;
wire \mreg/_00620_ ;
wire \mreg/_00621_ ;
wire \mreg/_00622_ ;
wire \mreg/_00623_ ;
wire \mreg/_00624_ ;
wire \mreg/_00625_ ;
wire \mreg/_00626_ ;
wire \mreg/_00627_ ;
wire \mreg/_00628_ ;
wire \mreg/_00629_ ;
wire \mreg/_00630_ ;
wire \mreg/_00631_ ;
wire \mreg/_00632_ ;
wire \mreg/_00633_ ;
wire \mreg/_00634_ ;
wire \mreg/_00635_ ;
wire \mreg/_00636_ ;
wire \mreg/_00637_ ;
wire \mreg/_00638_ ;
wire \mreg/_00639_ ;
wire \mreg/_00640_ ;
wire \mreg/_00641_ ;
wire \mreg/_00642_ ;
wire \mreg/_00643_ ;
wire \mreg/_00644_ ;
wire \mreg/_00645_ ;
wire \mreg/_00646_ ;
wire \mreg/_00647_ ;
wire \mreg/_00648_ ;
wire \mreg/_00649_ ;
wire \mreg/_00650_ ;
wire \mreg/_00651_ ;
wire \mreg/_00652_ ;
wire \mreg/_00653_ ;
wire \mreg/_00654_ ;
wire \mreg/_00655_ ;
wire \mreg/_00656_ ;
wire \mreg/_00657_ ;
wire \mreg/_00658_ ;
wire \mreg/_00659_ ;
wire \mreg/_00660_ ;
wire \mreg/_00661_ ;
wire \mreg/_00662_ ;
wire \mreg/_00663_ ;
wire \mreg/_00664_ ;
wire \mreg/_00665_ ;
wire \mreg/_00666_ ;
wire \mreg/_00667_ ;
wire \mreg/_00668_ ;
wire \mreg/_00669_ ;
wire \mreg/_00670_ ;
wire \mreg/_00671_ ;
wire \mreg/_00672_ ;
wire \mreg/_00673_ ;
wire \mreg/_00674_ ;
wire \mreg/_00675_ ;
wire \mreg/_00676_ ;
wire \mreg/_00677_ ;
wire \mreg/_00678_ ;
wire \mreg/_00679_ ;
wire \mreg/_00680_ ;
wire \mreg/_00681_ ;
wire \mreg/_00682_ ;
wire \mreg/_00683_ ;
wire \mreg/_00684_ ;
wire \mreg/_00685_ ;
wire \mreg/_00686_ ;
wire \mreg/_00687_ ;
wire \mreg/_00688_ ;
wire \mreg/_00689_ ;
wire \mreg/_00690_ ;
wire \mreg/_00691_ ;
wire \mreg/_00692_ ;
wire \mreg/_00693_ ;
wire \mreg/_00694_ ;
wire \mreg/_00695_ ;
wire \mreg/_00696_ ;
wire \mreg/_00697_ ;
wire \mreg/_00698_ ;
wire \mreg/_00699_ ;
wire \mreg/_00700_ ;
wire \mreg/_00701_ ;
wire \mreg/_00702_ ;
wire \mreg/_00703_ ;
wire \mreg/_00704_ ;
wire \mreg/_00705_ ;
wire \mreg/_00706_ ;
wire \mreg/_00707_ ;
wire \mreg/_00708_ ;
wire \mreg/_00709_ ;
wire \mreg/_00710_ ;
wire \mreg/_00711_ ;
wire \mreg/_00712_ ;
wire \mreg/_00713_ ;
wire \mreg/_00714_ ;
wire \mreg/_00715_ ;
wire \mreg/_00716_ ;
wire \mreg/_00717_ ;
wire \mreg/_00718_ ;
wire \mreg/_00719_ ;
wire \mreg/_00720_ ;
wire \mreg/_00721_ ;
wire \mreg/_00722_ ;
wire \mreg/_00723_ ;
wire \mreg/_00724_ ;
wire \mreg/_00725_ ;
wire \mreg/_00726_ ;
wire \mreg/_00727_ ;
wire \mreg/_00728_ ;
wire \mreg/_00729_ ;
wire \mreg/_00730_ ;
wire \mreg/_00731_ ;
wire \mreg/_00732_ ;
wire \mreg/_00733_ ;
wire \mreg/_00734_ ;
wire \mreg/_00735_ ;
wire \mreg/_00736_ ;
wire \mreg/_00737_ ;
wire \mreg/_00738_ ;
wire \mreg/_00739_ ;
wire \mreg/_00740_ ;
wire \mreg/_00741_ ;
wire \mreg/_00742_ ;
wire \mreg/_00743_ ;
wire \mreg/_00744_ ;
wire \mreg/_00745_ ;
wire \mreg/_00746_ ;
wire \mreg/_00747_ ;
wire \mreg/_00748_ ;
wire \mreg/_00749_ ;
wire \mreg/_00750_ ;
wire \mreg/_00751_ ;
wire \mreg/_00752_ ;
wire \mreg/_00753_ ;
wire \mreg/_00754_ ;
wire \mreg/_00755_ ;
wire \mreg/_00756_ ;
wire \mreg/_00757_ ;
wire \mreg/_00758_ ;
wire \mreg/_00759_ ;
wire \mreg/_00760_ ;
wire \mreg/_00761_ ;
wire \mreg/_00762_ ;
wire \mreg/_00763_ ;
wire \mreg/_00764_ ;
wire \mreg/_00765_ ;
wire \mreg/_00766_ ;
wire \mreg/_00767_ ;
wire \mreg/_00768_ ;
wire \mreg/_00769_ ;
wire \mreg/_00770_ ;
wire \mreg/_00771_ ;
wire \mreg/_00772_ ;
wire \mreg/_00773_ ;
wire \mreg/_00774_ ;
wire \mreg/_00775_ ;
wire \mreg/_00776_ ;
wire \mreg/_00777_ ;
wire \mreg/_00778_ ;
wire \mreg/_00779_ ;
wire \mreg/_00780_ ;
wire \mreg/_00781_ ;
wire \mreg/_00782_ ;
wire \mreg/_00783_ ;
wire \mreg/_00784_ ;
wire \mreg/_00785_ ;
wire \mreg/_00786_ ;
wire \mreg/_00787_ ;
wire \mreg/_00788_ ;
wire \mreg/_00789_ ;
wire \mreg/_00790_ ;
wire \mreg/_00791_ ;
wire \mreg/_00792_ ;
wire \mreg/_00793_ ;
wire \mreg/_00794_ ;
wire \mreg/_00795_ ;
wire \mreg/_00796_ ;
wire \mreg/_00797_ ;
wire \mreg/_00798_ ;
wire \mreg/_00799_ ;
wire \mreg/_00800_ ;
wire \mreg/_00801_ ;
wire \mreg/_00802_ ;
wire \mreg/_00803_ ;
wire \mreg/_00804_ ;
wire \mreg/_00805_ ;
wire \mreg/_00806_ ;
wire \mreg/_00807_ ;
wire \mreg/_00808_ ;
wire \mreg/_00809_ ;
wire \mreg/_00810_ ;
wire \mreg/_00811_ ;
wire \mreg/_00812_ ;
wire \mreg/_00813_ ;
wire \mreg/_00814_ ;
wire \mreg/_00815_ ;
wire \mreg/_00816_ ;
wire \mreg/_00817_ ;
wire \mreg/_00818_ ;
wire \mreg/_00819_ ;
wire \mreg/_00820_ ;
wire \mreg/_00821_ ;
wire \mreg/_00822_ ;
wire \mreg/_00823_ ;
wire \mreg/_00824_ ;
wire \mreg/_00825_ ;
wire \mreg/_00826_ ;
wire \mreg/_00827_ ;
wire \mreg/_00828_ ;
wire \mreg/_00829_ ;
wire \mreg/_00830_ ;
wire \mreg/_00831_ ;
wire \mreg/_00832_ ;
wire \mreg/_00833_ ;
wire \mreg/_00834_ ;
wire \mreg/_00835_ ;
wire \mreg/_00836_ ;
wire \mreg/_00837_ ;
wire \mreg/_00838_ ;
wire \mreg/_00839_ ;
wire \mreg/_00840_ ;
wire \mreg/_00841_ ;
wire \mreg/_00842_ ;
wire \mreg/_00843_ ;
wire \mreg/_00844_ ;
wire \mreg/_00845_ ;
wire \mreg/_00846_ ;
wire \mreg/_00847_ ;
wire \mreg/_00848_ ;
wire \mreg/_00849_ ;
wire \mreg/_00850_ ;
wire \mreg/_00851_ ;
wire \mreg/_00852_ ;
wire \mreg/_00853_ ;
wire \mreg/_00854_ ;
wire \mreg/_00855_ ;
wire \mreg/_00856_ ;
wire \mreg/_00857_ ;
wire \mreg/_00858_ ;
wire \mreg/_00859_ ;
wire \mreg/_00860_ ;
wire \mreg/_00861_ ;
wire \mreg/_00862_ ;
wire \mreg/_00863_ ;
wire \mreg/_00864_ ;
wire \mreg/_00865_ ;
wire \mreg/_00866_ ;
wire \mreg/_00867_ ;
wire \mreg/_00868_ ;
wire \mreg/_00869_ ;
wire \mreg/_00870_ ;
wire \mreg/_00871_ ;
wire \mreg/_00872_ ;
wire \mreg/_00873_ ;
wire \mreg/_00874_ ;
wire \mreg/_00875_ ;
wire \mreg/_00876_ ;
wire \mreg/_00877_ ;
wire \mreg/_00878_ ;
wire \mreg/_00879_ ;
wire \mreg/_00880_ ;
wire \mreg/_00881_ ;
wire \mreg/_00882_ ;
wire \mreg/_00883_ ;
wire \mreg/_00884_ ;
wire \mreg/_00885_ ;
wire \mreg/_00886_ ;
wire \mreg/_00887_ ;
wire \mreg/_00888_ ;
wire \mreg/_00889_ ;
wire \mreg/_00890_ ;
wire \mreg/_00891_ ;
wire \mreg/_00892_ ;
wire \mreg/_00893_ ;
wire \mreg/_00894_ ;
wire \mreg/_00895_ ;
wire \mreg/_00896_ ;
wire \mreg/_00897_ ;
wire \mreg/_00898_ ;
wire \mreg/_00899_ ;
wire \mreg/_00900_ ;
wire \mreg/_00901_ ;
wire \mreg/_00902_ ;
wire \mreg/_00903_ ;
wire \mreg/_00904_ ;
wire \mreg/_00905_ ;
wire \mreg/_00906_ ;
wire \mreg/_00907_ ;
wire \mreg/_00908_ ;
wire \mreg/_00909_ ;
wire \mreg/_00910_ ;
wire \mreg/_00911_ ;
wire \mreg/_00912_ ;
wire \mreg/_00913_ ;
wire \mreg/_00914_ ;
wire \mreg/_00915_ ;
wire \mreg/_00916_ ;
wire \mreg/_00917_ ;
wire \mreg/_00918_ ;
wire \mreg/_00919_ ;
wire \mreg/_00920_ ;
wire \mreg/_00921_ ;
wire \mreg/_00922_ ;
wire \mreg/_00923_ ;
wire \mreg/_00924_ ;
wire \mreg/_00925_ ;
wire \mreg/_00926_ ;
wire \mreg/_00927_ ;
wire \mreg/_00928_ ;
wire \mreg/_00929_ ;
wire \mreg/_00930_ ;
wire \mreg/_00931_ ;
wire \mreg/_00932_ ;
wire \mreg/_00933_ ;
wire \mreg/_00934_ ;
wire \mreg/_00935_ ;
wire \mreg/_00936_ ;
wire \mreg/_00937_ ;
wire \mreg/_00938_ ;
wire \mreg/_00939_ ;
wire \mreg/_00940_ ;
wire \mreg/_00941_ ;
wire \mreg/_00942_ ;
wire \mreg/_00943_ ;
wire \mreg/_00944_ ;
wire \mreg/_00945_ ;
wire \mreg/_00946_ ;
wire \mreg/_00947_ ;
wire \mreg/_00948_ ;
wire \mreg/_00949_ ;
wire \mreg/_00950_ ;
wire \mreg/_00951_ ;
wire \mreg/_00952_ ;
wire \mreg/_00953_ ;
wire \mreg/_00954_ ;
wire \mreg/_00955_ ;
wire \mreg/_00956_ ;
wire \mreg/_00957_ ;
wire \mreg/_00958_ ;
wire \mreg/_00959_ ;
wire \mreg/_00960_ ;
wire \mreg/_00961_ ;
wire \mreg/_00962_ ;
wire \mreg/_00963_ ;
wire \mreg/_00964_ ;
wire \mreg/_00965_ ;
wire \mreg/_00966_ ;
wire \mreg/_00967_ ;
wire \mreg/_00968_ ;
wire \mreg/_00969_ ;
wire \mreg/_00970_ ;
wire \mreg/_00971_ ;
wire \mreg/_00972_ ;
wire \mreg/_00973_ ;
wire \mreg/_00974_ ;
wire \mreg/_00975_ ;
wire \mreg/_00976_ ;
wire \mreg/_00977_ ;
wire \mreg/_00978_ ;
wire \mreg/_00979_ ;
wire \mreg/_00980_ ;
wire \mreg/_00981_ ;
wire \mreg/_00982_ ;
wire \mreg/_00983_ ;
wire \mreg/_00984_ ;
wire \mreg/_00985_ ;
wire \mreg/_00986_ ;
wire \mreg/_00987_ ;
wire \mreg/_00988_ ;
wire \mreg/_00989_ ;
wire \mreg/_00990_ ;
wire \mreg/_00991_ ;
wire \mreg/_00992_ ;
wire \mreg/_00993_ ;
wire \mreg/_00994_ ;
wire \mreg/_00995_ ;
wire \mreg/_00996_ ;
wire \mreg/_00997_ ;
wire \mreg/_00998_ ;
wire \mreg/_00999_ ;
wire \mreg/_01000_ ;
wire \mreg/_01001_ ;
wire \mreg/_01002_ ;
wire \mreg/_01003_ ;
wire \mreg/_01004_ ;
wire \mreg/_01005_ ;
wire \mreg/_01006_ ;
wire \mreg/_01007_ ;
wire \mreg/_01008_ ;
wire \mreg/_01009_ ;
wire \mreg/_01010_ ;
wire \mreg/_01011_ ;
wire \mreg/_01012_ ;
wire \mreg/_01013_ ;
wire \mreg/_01014_ ;
wire \mreg/_01015_ ;
wire \mreg/_01016_ ;
wire \mreg/_01017_ ;
wire \mreg/_01018_ ;
wire \mreg/_01019_ ;
wire \mreg/_01020_ ;
wire \mreg/_01021_ ;
wire \mreg/_01022_ ;
wire \mreg/_01023_ ;
wire \mreg/_01024_ ;
wire \mreg/_01025_ ;
wire \mreg/_01026_ ;
wire \mreg/_01027_ ;
wire \mreg/_01028_ ;
wire \mreg/_01029_ ;
wire \mreg/_01030_ ;
wire \mreg/_01031_ ;
wire \mreg/_01032_ ;
wire \mreg/_01033_ ;
wire \mreg/_01034_ ;
wire \mreg/_01035_ ;
wire \mreg/_01036_ ;
wire \mreg/_01037_ ;
wire \mreg/_01038_ ;
wire \mreg/_01039_ ;
wire \mreg/_01040_ ;
wire \mreg/_01041_ ;
wire \mreg/_01042_ ;
wire \mreg/_01043_ ;
wire \mreg/_01044_ ;
wire \mreg/_01045_ ;
wire \mreg/_01046_ ;
wire \mreg/_01047_ ;
wire \mreg/_01048_ ;
wire \mreg/_01049_ ;
wire \mreg/_01050_ ;
wire \mreg/_01051_ ;
wire \mreg/_01052_ ;
wire \mreg/_01053_ ;
wire \mreg/_01054_ ;
wire \mreg/_01055_ ;
wire \mreg/_01056_ ;
wire \mreg/_01057_ ;
wire \mreg/_01058_ ;
wire \mreg/_01059_ ;
wire \mreg/_01060_ ;
wire \mreg/_01061_ ;
wire \mreg/_01062_ ;
wire \mreg/_01063_ ;
wire \mreg/_01064_ ;
wire \mreg/_01065_ ;
wire \mreg/_01066_ ;
wire \mreg/_01067_ ;
wire \mreg/_01068_ ;
wire \mreg/_01069_ ;
wire \mreg/_01070_ ;
wire \mreg/_01071_ ;
wire \mreg/_01072_ ;
wire \mreg/_01073_ ;
wire \mreg/_01074_ ;
wire \mreg/_01075_ ;
wire \mreg/_01076_ ;
wire \mreg/_01077_ ;
wire \mreg/_01078_ ;
wire \mreg/_01079_ ;
wire \mreg/_01080_ ;
wire \mreg/_01081_ ;
wire \mreg/_01082_ ;
wire \mreg/_01083_ ;
wire \mreg/_01084_ ;
wire \mreg/_01085_ ;
wire \mreg/_01086_ ;
wire \mreg/_01087_ ;
wire \mreg/_01088_ ;
wire \mreg/_01089_ ;
wire \mreg/_01090_ ;
wire \mreg/_01091_ ;
wire \mreg/_01092_ ;
wire \mreg/_01093_ ;
wire \mreg/_01094_ ;
wire \mreg/_01095_ ;
wire \mreg/_01096_ ;
wire \mreg/_01097_ ;
wire \mreg/_01098_ ;
wire \mreg/_01099_ ;
wire \mreg/_01100_ ;
wire \mreg/_01101_ ;
wire \mreg/_01102_ ;
wire \mreg/_01103_ ;
wire \mreg/_01104_ ;
wire \mreg/_01105_ ;
wire \mreg/_01106_ ;
wire \mreg/_01107_ ;
wire \mreg/_01108_ ;
wire \mreg/_01109_ ;
wire \mreg/_01110_ ;
wire \mreg/_01111_ ;
wire \mreg/_01112_ ;
wire \mreg/_01113_ ;
wire \mreg/_01114_ ;
wire \mreg/_01115_ ;
wire \mreg/_01116_ ;
wire \mreg/_01117_ ;
wire \mreg/_01118_ ;
wire \mreg/_01119_ ;
wire \mreg/_01120_ ;
wire \mreg/_01121_ ;
wire \mreg/_01122_ ;
wire \mreg/_01123_ ;
wire \mreg/_01124_ ;
wire \mreg/_01125_ ;
wire \mreg/_01126_ ;
wire \mreg/_01127_ ;
wire \mreg/_01128_ ;
wire \mreg/_01129_ ;
wire \mreg/_01130_ ;
wire \mreg/_01131_ ;
wire \mreg/_01132_ ;
wire \mreg/_01133_ ;
wire \mreg/_01134_ ;
wire \mreg/_01135_ ;
wire \mreg/_01136_ ;
wire \mreg/_01137_ ;
wire \mreg/_01138_ ;
wire \mreg/_01139_ ;
wire \mreg/_01140_ ;
wire \mreg/_01141_ ;
wire \mreg/_01142_ ;
wire \mreg/_01143_ ;
wire \mreg/_01144_ ;
wire \mreg/_01145_ ;
wire \mreg/_01146_ ;
wire \mreg/_01147_ ;
wire \mreg/_01148_ ;
wire \mreg/_01149_ ;
wire \mreg/_01150_ ;
wire \mreg/_01151_ ;
wire \mreg/_01152_ ;
wire \mreg/_01153_ ;
wire \mreg/_01154_ ;
wire \mreg/_01155_ ;
wire \mreg/_01156_ ;
wire \mreg/_01157_ ;
wire \mreg/_01158_ ;
wire \mreg/_01159_ ;
wire \mreg/_01160_ ;
wire \mreg/_01161_ ;
wire \mreg/_01162_ ;
wire \mreg/_01163_ ;
wire \mreg/_01164_ ;
wire \mreg/_01165_ ;
wire \mreg/_01166_ ;
wire \mreg/_01167_ ;
wire \mreg/_01168_ ;
wire \mreg/_01169_ ;
wire \mreg/_01170_ ;
wire \mreg/_01171_ ;
wire \mreg/_01172_ ;
wire \mreg/_01173_ ;
wire \mreg/_01174_ ;
wire \mreg/_01175_ ;
wire \mreg/_01176_ ;
wire \mreg/_01177_ ;
wire \mreg/_01178_ ;
wire \mreg/_01179_ ;
wire \mreg/_01180_ ;
wire \mreg/_01181_ ;
wire \mreg/_01182_ ;
wire \mreg/_01183_ ;
wire \mreg/_01184_ ;
wire \mreg/_01185_ ;
wire \mreg/_01186_ ;
wire \mreg/_01187_ ;
wire \mreg/_01188_ ;
wire \mreg/_01189_ ;
wire \mreg/_01190_ ;
wire \mreg/_01191_ ;
wire \mreg/_01192_ ;
wire \mreg/_01193_ ;
wire \mreg/_01194_ ;
wire \mreg/_01195_ ;
wire \mreg/_01196_ ;
wire \mreg/_01197_ ;
wire \mreg/_01198_ ;
wire \mreg/_01199_ ;
wire \mreg/_01200_ ;
wire \mreg/_01201_ ;
wire \mreg/_01202_ ;
wire \mreg/_01203_ ;
wire \mreg/_01204_ ;
wire \mreg/_01205_ ;
wire \mreg/_01206_ ;
wire \mreg/_01207_ ;
wire \mreg/_01208_ ;
wire \mreg/_01209_ ;
wire \mreg/_01210_ ;
wire \mreg/_01211_ ;
wire \mreg/_01212_ ;
wire \mreg/_01213_ ;
wire \mreg/_01214_ ;
wire \mreg/_01215_ ;
wire \mreg/_01216_ ;
wire \mreg/_01217_ ;
wire \mreg/_01218_ ;
wire \mreg/_01219_ ;
wire \mreg/_01220_ ;
wire \mreg/_01221_ ;
wire \mreg/_01222_ ;
wire \mreg/_01223_ ;
wire \mreg/_01224_ ;
wire \mreg/_01225_ ;
wire \mreg/_01226_ ;
wire \mreg/_01227_ ;
wire \mreg/_01228_ ;
wire \mreg/_01229_ ;
wire \mreg/_01230_ ;
wire \mreg/_01231_ ;
wire \mreg/_01232_ ;
wire \mreg/_01233_ ;
wire \mreg/_01234_ ;
wire \mreg/_01235_ ;
wire \mreg/_01236_ ;
wire \mreg/_01237_ ;
wire \mreg/_01238_ ;
wire \mreg/_01239_ ;
wire \mreg/_01240_ ;
wire \mreg/_01241_ ;
wire \mreg/_01242_ ;
wire \mreg/_01243_ ;
wire \mreg/_01244_ ;
wire \mreg/_01245_ ;
wire \mreg/_01246_ ;
wire \mreg/_01247_ ;
wire \mreg/_01248_ ;
wire \mreg/_01249_ ;
wire \mreg/_01250_ ;
wire \mreg/_01251_ ;
wire \mreg/_01252_ ;
wire \mreg/_01253_ ;
wire \mreg/_01254_ ;
wire \mreg/_01255_ ;
wire \mreg/_01256_ ;
wire \mreg/_01257_ ;
wire \mreg/_01258_ ;
wire \mreg/_01259_ ;
wire \mreg/_01260_ ;
wire \mreg/_01261_ ;
wire \mreg/_01262_ ;
wire \mreg/_01263_ ;
wire \mreg/_01264_ ;
wire \mreg/_01265_ ;
wire \mreg/_01266_ ;
wire \mreg/_01267_ ;
wire \mreg/_01268_ ;
wire \mreg/_01269_ ;
wire \mreg/_01270_ ;
wire \mreg/_01271_ ;
wire \mreg/_01272_ ;
wire \mreg/_01273_ ;
wire \mreg/_01274_ ;
wire \mreg/_01275_ ;
wire \mreg/_01276_ ;
wire \mreg/_01277_ ;
wire \mreg/_01278_ ;
wire \mreg/_01279_ ;
wire \mreg/_01280_ ;
wire \mreg/_01281_ ;
wire \mreg/_01282_ ;
wire \mreg/_01283_ ;
wire \mreg/_01284_ ;
wire \mreg/_01285_ ;
wire \mreg/_01286_ ;
wire \mreg/_01287_ ;
wire \mreg/_01288_ ;
wire \mreg/_01289_ ;
wire \mreg/_01290_ ;
wire \mreg/_01291_ ;
wire \mreg/_01292_ ;
wire \mreg/_01293_ ;
wire \mreg/_01294_ ;
wire \mreg/_01295_ ;
wire \mreg/_01296_ ;
wire \mreg/_01297_ ;
wire \mreg/_01298_ ;
wire \mreg/_01299_ ;
wire \mreg/_01300_ ;
wire \mreg/_01301_ ;
wire \mreg/_01302_ ;
wire \mreg/_01303_ ;
wire \mreg/_01304_ ;
wire \mreg/_01305_ ;
wire \mreg/_01306_ ;
wire \mreg/_01307_ ;
wire \mreg/_01308_ ;
wire \mreg/_01309_ ;
wire \mreg/_01310_ ;
wire \mreg/_01311_ ;
wire \mreg/_01312_ ;
wire \mreg/_01313_ ;
wire \mreg/_01314_ ;
wire \mreg/_01315_ ;
wire \mreg/_01316_ ;
wire \mreg/_01317_ ;
wire \mreg/_01318_ ;
wire \mreg/_01319_ ;
wire \mreg/_01320_ ;
wire \mreg/_01321_ ;
wire \mreg/_01322_ ;
wire \mreg/_01323_ ;
wire \mreg/_01324_ ;
wire \mreg/_01325_ ;
wire \mreg/_01326_ ;
wire \mreg/_01327_ ;
wire \mreg/_01328_ ;
wire \mreg/_01329_ ;
wire \mreg/_01330_ ;
wire \mreg/_01331_ ;
wire \mreg/_01332_ ;
wire \mreg/_01333_ ;
wire \mreg/_01334_ ;
wire \mreg/_01335_ ;
wire \mreg/_01336_ ;
wire \mreg/_01337_ ;
wire \mreg/_01338_ ;
wire \mreg/_01339_ ;
wire \mreg/_01340_ ;
wire \mreg/_01341_ ;
wire \mreg/_01342_ ;
wire \mreg/_01343_ ;
wire \mreg/_01344_ ;
wire \mreg/_01345_ ;
wire \mreg/_01346_ ;
wire \mreg/_01347_ ;
wire \mreg/_01348_ ;
wire \mreg/_01349_ ;
wire \mreg/_01350_ ;
wire \mreg/_01351_ ;
wire \mreg/_01352_ ;
wire \mreg/_01353_ ;
wire \mreg/_01354_ ;
wire \mreg/_01355_ ;
wire \mreg/_01356_ ;
wire \mreg/_01357_ ;
wire \mreg/_01358_ ;
wire \mreg/_01359_ ;
wire \mreg/_01360_ ;
wire \mreg/_01361_ ;
wire \mreg/_01362_ ;
wire \mreg/_01363_ ;
wire \mreg/_01364_ ;
wire \mreg/_01365_ ;
wire \mreg/_01366_ ;
wire \mreg/_01367_ ;
wire \mreg/_01368_ ;
wire \mreg/_01369_ ;
wire \mreg/_01370_ ;
wire \mreg/_01371_ ;
wire \mreg/_01372_ ;
wire \mreg/_01373_ ;
wire \mreg/_01374_ ;
wire \mreg/_01375_ ;
wire \mreg/_01376_ ;
wire \mreg/_01377_ ;
wire \mreg/_01378_ ;
wire \mreg/_01379_ ;
wire \mreg/_01380_ ;
wire \mreg/_01381_ ;
wire \mreg/_01382_ ;
wire \mreg/_01383_ ;
wire \mreg/_01384_ ;
wire \mreg/_01385_ ;
wire \mreg/_01386_ ;
wire \mreg/_01387_ ;
wire \mreg/_01388_ ;
wire \mreg/_01389_ ;
wire \mreg/_01390_ ;
wire \mreg/_01391_ ;
wire \mreg/_01392_ ;
wire \mreg/_01393_ ;
wire \mreg/_01394_ ;
wire \mreg/_01395_ ;
wire \mreg/_01396_ ;
wire \mreg/_01397_ ;
wire \mreg/_01398_ ;
wire \mreg/_01399_ ;
wire \mreg/_01400_ ;
wire \mreg/_01401_ ;
wire \mreg/_01402_ ;
wire \mreg/_01403_ ;
wire \mreg/_01404_ ;
wire \mreg/_01405_ ;
wire \mreg/_01406_ ;
wire \mreg/_01407_ ;
wire \mreg/_01408_ ;
wire \mreg/_01409_ ;
wire \mreg/_01410_ ;
wire \mreg/_01411_ ;
wire \mreg/_01412_ ;
wire \mreg/_01413_ ;
wire \mreg/_01414_ ;
wire \mreg/_01415_ ;
wire \mreg/_01416_ ;
wire \mreg/_01417_ ;
wire \mreg/_01418_ ;
wire \mreg/_01419_ ;
wire \mreg/_01420_ ;
wire \mreg/_01421_ ;
wire \mreg/_01422_ ;
wire \mreg/_01423_ ;
wire \mreg/_01424_ ;
wire \mreg/_01425_ ;
wire \mreg/_01426_ ;
wire \mreg/_01427_ ;
wire \mreg/_01428_ ;
wire \mreg/_01429_ ;
wire \mreg/_01430_ ;
wire \mreg/_01431_ ;
wire \mreg/_01432_ ;
wire \mreg/_01433_ ;
wire \mreg/_01434_ ;
wire \mreg/_01435_ ;
wire \mreg/_01436_ ;
wire \mreg/_01437_ ;
wire \mreg/_01438_ ;
wire \mreg/_01439_ ;
wire \mreg/_01440_ ;
wire \mreg/_01441_ ;
wire \mreg/_01442_ ;
wire \mreg/_01443_ ;
wire \mreg/_01444_ ;
wire \mreg/_01445_ ;
wire \mreg/_01446_ ;
wire \mreg/_01447_ ;
wire \mreg/_01448_ ;
wire \mreg/_01449_ ;
wire \mreg/_01450_ ;
wire \mreg/_01451_ ;
wire \mreg/_01452_ ;
wire \mreg/_01453_ ;
wire \mreg/_01454_ ;
wire \mreg/_01455_ ;
wire \mreg/_01456_ ;
wire \mreg/_01457_ ;
wire \mreg/_01458_ ;
wire \mreg/_01459_ ;
wire \mreg/_01460_ ;
wire \mreg/_01461_ ;
wire \mreg/_01462_ ;
wire \mreg/_01463_ ;
wire \mreg/_01464_ ;
wire \mreg/_01465_ ;
wire \mreg/_01466_ ;
wire \mreg/_01467_ ;
wire \mreg/_01468_ ;
wire \mreg/_01469_ ;
wire \mreg/_01470_ ;
wire \mreg/_01471_ ;
wire \mreg/_01472_ ;
wire \mreg/_01473_ ;
wire \mreg/_01474_ ;
wire \mreg/_01475_ ;
wire \mreg/_01476_ ;
wire \mreg/_01477_ ;
wire \mreg/_01478_ ;
wire \mreg/_01479_ ;
wire \mreg/_01480_ ;
wire \mreg/_01481_ ;
wire \mreg/_01482_ ;
wire \mreg/_01483_ ;
wire \mreg/_01484_ ;
wire \mreg/_01485_ ;
wire \mreg/_01486_ ;
wire \mreg/_01487_ ;
wire \mreg/_01488_ ;
wire \mreg/_01489_ ;
wire \mreg/_01490_ ;
wire \mreg/_01491_ ;
wire \mreg/_01492_ ;
wire \mreg/_01493_ ;
wire \mreg/_01494_ ;
wire \mreg/_01495_ ;
wire \mreg/_01496_ ;
wire \mreg/_01497_ ;
wire \mreg/_01498_ ;
wire \mreg/_01499_ ;
wire \mreg/_01500_ ;
wire \mreg/_01501_ ;
wire \mreg/_01502_ ;
wire \mreg/_01503_ ;
wire \mreg/_01504_ ;
wire \mreg/_01505_ ;
wire \mreg/_01506_ ;
wire \mreg/_01507_ ;
wire \mreg/_01508_ ;
wire \mreg/_01509_ ;
wire \mreg/_01510_ ;
wire \mreg/_01511_ ;
wire \mreg/_01512_ ;
wire \mreg/_01513_ ;
wire \mreg/_01514_ ;
wire \mreg/_01515_ ;
wire \mreg/_01516_ ;
wire \mreg/_01517_ ;
wire \mreg/_01518_ ;
wire \mreg/_01519_ ;
wire \mreg/_01520_ ;
wire \mreg/_01521_ ;
wire \mreg/_01522_ ;
wire \mreg/_01523_ ;
wire \mreg/_01524_ ;
wire \mreg/_01525_ ;
wire \mreg/_01526_ ;
wire \mreg/_01527_ ;
wire \mreg/_01528_ ;
wire \mreg/_01529_ ;
wire \mreg/_01530_ ;
wire \mreg/_01531_ ;
wire \mreg/_01532_ ;
wire \mreg/_01533_ ;
wire \mreg/_01534_ ;
wire \mreg/_01535_ ;
wire \mreg/_01536_ ;
wire \mreg/_01537_ ;
wire \mreg/_01538_ ;
wire \mreg/_01539_ ;
wire \mreg/_01540_ ;
wire \mreg/_01541_ ;
wire \mreg/_01542_ ;
wire \mreg/_01543_ ;
wire \mreg/_01544_ ;
wire \mreg/_01545_ ;
wire \mreg/_01546_ ;
wire \mreg/_01547_ ;
wire \mreg/_01548_ ;
wire \mreg/_01549_ ;
wire \mreg/_01550_ ;
wire \mreg/_01551_ ;
wire \mreg/_01552_ ;
wire \mreg/_01553_ ;
wire \mreg/_01554_ ;
wire \mreg/_01555_ ;
wire \mreg/_01556_ ;
wire \mreg/_01557_ ;
wire \mreg/_01558_ ;
wire \mreg/_01559_ ;
wire \mreg/_01560_ ;
wire \mreg/_01561_ ;
wire \mreg/_01562_ ;
wire \mreg/_01563_ ;
wire \mreg/_01564_ ;
wire \mreg/_01565_ ;
wire \mreg/_01566_ ;
wire \mreg/_01567_ ;
wire \mreg/_01568_ ;
wire \mreg/_01569_ ;
wire \mreg/_01570_ ;
wire \mreg/_01571_ ;
wire \mreg/_01572_ ;
wire \mreg/_01573_ ;
wire \mreg/_01574_ ;
wire \mreg/_01575_ ;
wire \mreg/_01576_ ;
wire \mreg/_01577_ ;
wire \mreg/_01578_ ;
wire \mreg/_01579_ ;
wire \mreg/_01580_ ;
wire \mreg/_01581_ ;
wire \mreg/_01582_ ;
wire \mreg/_01583_ ;
wire \mreg/_01584_ ;
wire \mreg/_01585_ ;
wire \mreg/_01586_ ;
wire \mreg/_01587_ ;
wire \mreg/_01588_ ;
wire \mreg/_01589_ ;
wire \mreg/_01590_ ;
wire \mreg/_01591_ ;
wire \mreg/_01592_ ;
wire \mreg/_01593_ ;
wire \mreg/_01594_ ;
wire \mreg/_01595_ ;
wire \mreg/_01596_ ;
wire \mreg/_01597_ ;
wire \mreg/_01598_ ;
wire \mreg/_01599_ ;
wire \mreg/_01600_ ;
wire \mreg/_01601_ ;
wire \mreg/_01602_ ;
wire \mreg/_01603_ ;
wire \mreg/_01604_ ;
wire \mreg/_01605_ ;
wire \mreg/_01606_ ;
wire \mreg/_01607_ ;
wire \mreg/_01608_ ;
wire \mreg/_01609_ ;
wire \mreg/_01610_ ;
wire \mreg/_01611_ ;
wire \mreg/_01612_ ;
wire \mreg/_01613_ ;
wire \mreg/_01614_ ;
wire \mreg/_01615_ ;
wire \mreg/_01616_ ;
wire \mreg/_01617_ ;
wire \mreg/_01618_ ;
wire \mreg/_01619_ ;
wire \mreg/_01620_ ;
wire \mreg/_01621_ ;
wire \mreg/_01622_ ;
wire \mreg/_01623_ ;
wire \mreg/_01624_ ;
wire \mreg/_01625_ ;
wire \mreg/_01626_ ;
wire \mreg/_01627_ ;
wire \mreg/_01628_ ;
wire \mreg/_01629_ ;
wire \mreg/_01630_ ;
wire \mreg/_01631_ ;
wire \mreg/_01632_ ;
wire \mreg/_01633_ ;
wire \mreg/_01634_ ;
wire \mreg/_01635_ ;
wire \mreg/_01636_ ;
wire \mreg/_01637_ ;
wire \mreg/_01638_ ;
wire \mreg/_01639_ ;
wire \mreg/_01640_ ;
wire \mreg/_01641_ ;
wire \mreg/_01642_ ;
wire \mreg/_01643_ ;
wire \mreg/_01644_ ;
wire \mreg/_01645_ ;
wire \mreg/_01646_ ;
wire \mreg/_01647_ ;
wire \mreg/_01648_ ;
wire \mreg/_01649_ ;
wire \mreg/_01650_ ;
wire \mreg/_01651_ ;
wire \mreg/_01652_ ;
wire \mreg/_01653_ ;
wire \mreg/_01654_ ;
wire \mreg/_01655_ ;
wire \mreg/_01656_ ;
wire \mreg/_01657_ ;
wire \mreg/_01658_ ;
wire \mreg/_01659_ ;
wire \mreg/_01660_ ;
wire \mreg/_01661_ ;
wire \mreg/_01662_ ;
wire \mreg/_01663_ ;
wire \mreg/_01664_ ;
wire \mreg/_01665_ ;
wire \mreg/_01666_ ;
wire \mreg/_01667_ ;
wire \mreg/_01668_ ;
wire \mreg/_01669_ ;
wire \mreg/_01670_ ;
wire \mreg/_01671_ ;
wire \mreg/_01672_ ;
wire \mreg/_01673_ ;
wire \mreg/_01674_ ;
wire \mreg/_01675_ ;
wire \mreg/_01676_ ;
wire \mreg/_01677_ ;
wire \mreg/_01678_ ;
wire \mreg/_01679_ ;
wire \mreg/_01680_ ;
wire \mreg/_01681_ ;
wire \mreg/_01682_ ;
wire \mreg/_01683_ ;
wire \mreg/_01684_ ;
wire \mreg/_01685_ ;
wire \mreg/_01686_ ;
wire \mreg/_01687_ ;
wire \mreg/_01688_ ;
wire \mreg/_01689_ ;
wire \mreg/_01690_ ;
wire \mreg/_01691_ ;
wire \mreg/_01692_ ;
wire \mreg/_01693_ ;
wire \mreg/_01694_ ;
wire \mreg/_01695_ ;
wire \mreg/_01696_ ;
wire \mreg/_01697_ ;
wire \mreg/_01698_ ;
wire \mreg/_01699_ ;
wire \mreg/_01700_ ;
wire \mreg/_01701_ ;
wire \mreg/_01702_ ;
wire \mreg/_01703_ ;
wire \mreg/_01704_ ;
wire \mreg/_01705_ ;
wire \mreg/_01706_ ;
wire \mreg/_01707_ ;
wire \mreg/_01708_ ;
wire \mreg/_01709_ ;
wire \mreg/_01710_ ;
wire \mreg/_01711_ ;
wire \mreg/_01712_ ;
wire \mreg/_01713_ ;
wire \mreg/_01714_ ;
wire \mreg/_01715_ ;
wire \mreg/_01716_ ;
wire \mreg/_01717_ ;
wire \mreg/_01718_ ;
wire \mreg/_01719_ ;
wire \mreg/_01720_ ;
wire \mreg/_01721_ ;
wire \mreg/_01722_ ;
wire \mreg/_01723_ ;
wire \mreg/_01724_ ;
wire \mreg/_01725_ ;
wire \mreg/_01726_ ;
wire \mreg/_01727_ ;
wire \mreg/_01728_ ;
wire \mreg/_01729_ ;
wire \mreg/_01730_ ;
wire \mreg/_01731_ ;
wire \mreg/_01732_ ;
wire \mreg/_01733_ ;
wire \mreg/_01734_ ;
wire \mreg/_01735_ ;
wire \mreg/_01736_ ;
wire \mreg/_01737_ ;
wire \mreg/_01738_ ;
wire \mreg/_01739_ ;
wire \mreg/_01740_ ;
wire \mreg/_01741_ ;
wire \mreg/_01742_ ;
wire \mreg/_01743_ ;
wire \mreg/_01744_ ;
wire \mreg/_01745_ ;
wire \mreg/_01746_ ;
wire \mreg/_01747_ ;
wire \mreg/_01748_ ;
wire \mreg/_01749_ ;
wire \mreg/_01750_ ;
wire \mreg/_01751_ ;
wire \mreg/_01752_ ;
wire \mreg/_01753_ ;
wire \mreg/_01754_ ;
wire \mreg/_01755_ ;
wire \mreg/_01756_ ;
wire \mreg/_01757_ ;
wire \mreg/_01758_ ;
wire \mreg/_01759_ ;
wire \mreg/_01760_ ;
wire \mreg/_01761_ ;
wire \mreg/_01762_ ;
wire \mreg/_01763_ ;
wire \mreg/_01764_ ;
wire \mreg/_01765_ ;
wire \mreg/_01766_ ;
wire \mreg/_01767_ ;
wire \mreg/_01768_ ;
wire \mreg/_01769_ ;
wire \mreg/_01770_ ;
wire \mreg/_01771_ ;
wire \mreg/_01772_ ;
wire \mreg/_01773_ ;
wire \mreg/_01774_ ;
wire \mreg/_01775_ ;
wire \mreg/_01776_ ;
wire \mreg/_01777_ ;
wire \mreg/_01778_ ;
wire \mreg/_01779_ ;
wire \mreg/_01780_ ;
wire \mreg/_01781_ ;
wire \mreg/_01782_ ;
wire \mreg/_01783_ ;
wire \mreg/_01784_ ;
wire \mreg/_01785_ ;
wire \mreg/_01786_ ;
wire \mreg/_01787_ ;
wire \mreg/_01788_ ;
wire \mreg/_01789_ ;
wire \mreg/_01790_ ;
wire \mreg/_01791_ ;
wire \mreg/_01792_ ;
wire \mreg/_01793_ ;
wire \mreg/_01794_ ;
wire \mreg/_01795_ ;
wire \mreg/_01796_ ;
wire \mreg/_01797_ ;
wire \mreg/_01798_ ;
wire \mreg/_01799_ ;
wire \mreg/_01800_ ;
wire \mreg/_01801_ ;
wire \mreg/_01802_ ;
wire \mreg/_01803_ ;
wire \mreg/_01804_ ;
wire \mreg/_01805_ ;
wire \mreg/_01806_ ;
wire \mreg/_01807_ ;
wire \mreg/_01808_ ;
wire \mreg/_01809_ ;
wire \mreg/_01810_ ;
wire \mreg/_01811_ ;
wire \mreg/_01812_ ;
wire \mreg/_01813_ ;
wire \mreg/_01814_ ;
wire \mreg/_01815_ ;
wire \mreg/_01816_ ;
wire \mreg/_01817_ ;
wire \mreg/_01818_ ;
wire \mreg/_01819_ ;
wire \mreg/_01820_ ;
wire \mreg/_01821_ ;
wire \mreg/_01822_ ;
wire \mreg/_01823_ ;
wire \mreg/_01824_ ;
wire \mreg/_01825_ ;
wire \mreg/_01826_ ;
wire \mreg/_01827_ ;
wire \mreg/_01828_ ;
wire \mreg/_01829_ ;
wire \mreg/_01830_ ;
wire \mreg/_01831_ ;
wire \mreg/_01832_ ;
wire \mreg/_01833_ ;
wire \mreg/_01834_ ;
wire \mreg/_01835_ ;
wire \mreg/_01836_ ;
wire \mreg/_01837_ ;
wire \mreg/_01838_ ;
wire \mreg/_01839_ ;
wire \mreg/_01840_ ;
wire \mreg/_01841_ ;
wire \mreg/_01842_ ;
wire \mreg/_01843_ ;
wire \mreg/_01844_ ;
wire \mreg/_01845_ ;
wire \mreg/_01846_ ;
wire \mreg/_01847_ ;
wire \mreg/_01848_ ;
wire \mreg/_01849_ ;
wire \mreg/_01850_ ;
wire \mreg/_01851_ ;
wire \mreg/_01852_ ;
wire \mreg/_01853_ ;
wire \mreg/_01854_ ;
wire \mreg/_01855_ ;
wire \mreg/_01856_ ;
wire \mreg/_01857_ ;
wire \mreg/_01858_ ;
wire \mreg/_01859_ ;
wire \mreg/_01860_ ;
wire \mreg/_01861_ ;
wire \mreg/_01862_ ;
wire \mreg/_01863_ ;
wire \mreg/_01864_ ;
wire \mreg/_01865_ ;
wire \mreg/_01866_ ;
wire \mreg/_01867_ ;
wire \mreg/_01868_ ;
wire \mreg/_01869_ ;
wire \mreg/_01870_ ;
wire \mreg/_01871_ ;
wire \mreg/_01872_ ;
wire \mreg/_01873_ ;
wire \mreg/_01874_ ;
wire \mreg/_01875_ ;
wire \mreg/_01876_ ;
wire \mreg/_01877_ ;
wire \mreg/_01878_ ;
wire \mreg/_01879_ ;
wire \mreg/_01880_ ;
wire \mreg/_01881_ ;
wire \mreg/_01882_ ;
wire \mreg/_01883_ ;
wire \mreg/_01884_ ;
wire \mreg/_01885_ ;
wire \mreg/_01886_ ;
wire \mreg/_01887_ ;
wire \mreg/_01888_ ;
wire \mreg/_01889_ ;
wire \mreg/_01890_ ;
wire \mreg/_01891_ ;
wire \mreg/_01892_ ;
wire \mreg/_01893_ ;
wire \mreg/_01894_ ;
wire \mreg/_01895_ ;
wire \mreg/_01896_ ;
wire \mreg/_01897_ ;
wire \mreg/_01898_ ;
wire \mreg/_01899_ ;
wire \mreg/_01900_ ;
wire \mreg/_01901_ ;
wire \mreg/_01902_ ;
wire \mreg/_01903_ ;
wire \mreg/_01904_ ;
wire \mreg/_01905_ ;
wire \mreg/_01906_ ;
wire \mreg/_01907_ ;
wire \mreg/_01908_ ;
wire \mreg/_01909_ ;
wire \mreg/_01910_ ;
wire \mreg/_01911_ ;
wire \mreg/_01912_ ;
wire \mreg/_01913_ ;
wire \mreg/_01914_ ;
wire \mreg/_01915_ ;
wire \mreg/_01916_ ;
wire \mreg/_01917_ ;
wire \mreg/_01918_ ;
wire \mreg/_01919_ ;
wire \mreg/_01920_ ;
wire \mreg/_01921_ ;
wire \mreg/_01922_ ;
wire \mreg/_01923_ ;
wire \mreg/_01924_ ;
wire \mreg/_01925_ ;
wire \mreg/_01926_ ;
wire \mreg/_01927_ ;
wire \mreg/_01928_ ;
wire \mreg/_01929_ ;
wire \mreg/_01930_ ;
wire \mreg/_01931_ ;
wire \mreg/_01932_ ;
wire \mreg/_01933_ ;
wire \mreg/_01934_ ;
wire \mreg/_01935_ ;
wire \mreg/_01936_ ;
wire \mreg/_01937_ ;
wire \mreg/_01938_ ;
wire \mreg/_01939_ ;
wire \mreg/_01940_ ;
wire \mreg/_01941_ ;
wire \mreg/_01942_ ;
wire \mreg/_01943_ ;
wire \mreg/_01944_ ;
wire \mreg/_01945_ ;
wire \mreg/_01946_ ;
wire \mreg/_01947_ ;
wire \mreg/_01948_ ;
wire \mreg/_01949_ ;
wire \mreg/_01950_ ;
wire \mreg/_01951_ ;
wire \mreg/_01952_ ;
wire \mreg/_01953_ ;
wire \mreg/_01954_ ;
wire \mreg/_01955_ ;
wire \mreg/_01956_ ;
wire \mreg/_01957_ ;
wire \mreg/_01958_ ;
wire \mreg/_01959_ ;
wire \mreg/_01960_ ;
wire \mreg/_01961_ ;
wire \mreg/_01962_ ;
wire \mreg/_01963_ ;
wire \mreg/_01964_ ;
wire \mreg/_01965_ ;
wire \mreg/_01966_ ;
wire \mreg/_01967_ ;
wire \mreg/_01968_ ;
wire \mreg/_01969_ ;
wire \mreg/_01970_ ;
wire \mreg/_01971_ ;
wire \mreg/_01972_ ;
wire \mreg/_01973_ ;
wire \mreg/_01974_ ;
wire \mreg/_01975_ ;
wire \mreg/_01976_ ;
wire \mreg/_01977_ ;
wire \mreg/_01978_ ;
wire \mreg/_01979_ ;
wire \mreg/_01980_ ;
wire \mreg/_01981_ ;
wire \mreg/_01982_ ;
wire \mreg/_01983_ ;
wire \mreg/_01984_ ;
wire \mreg/_01985_ ;
wire \mreg/_01986_ ;
wire \mreg/_01987_ ;
wire \mreg/_01988_ ;
wire \mreg/_01989_ ;
wire \mreg/_01990_ ;
wire \mreg/_01991_ ;
wire \mreg/_01992_ ;
wire \mreg/_01993_ ;
wire \mreg/_01994_ ;
wire \mreg/_01995_ ;
wire \mreg/_01996_ ;
wire \mreg/_01997_ ;
wire \mreg/_01998_ ;
wire \mreg/_01999_ ;
wire \mreg/_02000_ ;
wire \mreg/_02001_ ;
wire \mreg/_02002_ ;
wire \mreg/_02003_ ;
wire \mreg/_02004_ ;
wire \mreg/_02005_ ;
wire \mreg/_02006_ ;
wire \mreg/_02007_ ;
wire \mreg/_02008_ ;
wire \mreg/_02009_ ;
wire \mreg/_02010_ ;
wire \mreg/_02011_ ;
wire \mreg/_02012_ ;
wire \mreg/_02013_ ;
wire \mreg/_02014_ ;
wire \mreg/_02015_ ;
wire \mreg/_02016_ ;
wire \mreg/_02017_ ;
wire \mreg/_02018_ ;
wire \mreg/_02019_ ;
wire \mreg/_02020_ ;
wire \mreg/_02021_ ;
wire \mreg/_02022_ ;
wire \mreg/_02023_ ;
wire \mreg/_02024_ ;
wire \mreg/_02025_ ;
wire \mreg/_02026_ ;
wire \mreg/_02027_ ;
wire \mreg/_02028_ ;
wire \mreg/_02029_ ;
wire \mreg/_02030_ ;
wire \mreg/_02031_ ;
wire \mreg/_02032_ ;
wire \mreg/_02033_ ;
wire \mreg/_02034_ ;
wire \mreg/_02035_ ;
wire \mreg/_02036_ ;
wire \mreg/_02037_ ;
wire \mreg/_02038_ ;
wire \mreg/_02039_ ;
wire \mreg/_02040_ ;
wire \mreg/_02041_ ;
wire \mreg/_02042_ ;
wire \mreg/_02043_ ;
wire \mreg/_02044_ ;
wire \mreg/_02045_ ;
wire \mreg/_02046_ ;
wire \mreg/_02047_ ;
wire \mreg/_02048_ ;
wire \mreg/_02049_ ;
wire \mreg/_02050_ ;
wire \mreg/_02051_ ;
wire \mreg/_02052_ ;
wire \mreg/_02053_ ;
wire \mreg/_02054_ ;
wire \mreg/_02055_ ;
wire \mreg/_02056_ ;
wire \mreg/_02057_ ;
wire \mreg/_02058_ ;
wire \mreg/_02059_ ;
wire \mreg/_02060_ ;
wire \mreg/_02061_ ;
wire \mreg/_02062_ ;
wire \mreg/_02063_ ;
wire \mreg/_02064_ ;
wire \mreg/_02065_ ;
wire \mreg/_02066_ ;
wire \mreg/_02067_ ;
wire \mreg/_02068_ ;
wire \mreg/_02069_ ;
wire \mreg/_02070_ ;
wire \mreg/_02071_ ;
wire \mreg/_02072_ ;
wire \mreg/_02073_ ;
wire \mreg/_02074_ ;
wire \mreg/_02075_ ;
wire \mreg/_02076_ ;
wire \mreg/_02077_ ;
wire \mreg/_02078_ ;
wire \mreg/_02079_ ;
wire \mreg/_02080_ ;
wire \mreg/_02081_ ;
wire \mreg/_02082_ ;
wire \mreg/_02083_ ;
wire \mreg/_02084_ ;
wire \mreg/_02085_ ;
wire \mreg/_02086_ ;
wire \mreg/_02087_ ;
wire \mreg/_02088_ ;
wire \mreg/_02089_ ;
wire \mreg/_02090_ ;
wire \mreg/_02091_ ;
wire \mreg/_02092_ ;
wire \mreg/_02093_ ;
wire \mreg/_02094_ ;
wire \mreg/_02095_ ;
wire \mreg/_02096_ ;
wire \mreg/_02097_ ;
wire \mreg/_02098_ ;
wire \mreg/_02099_ ;
wire \mreg/_02100_ ;
wire \mreg/_02101_ ;
wire \mreg/_02102_ ;
wire \mreg/_02103_ ;
wire \mreg/_02104_ ;
wire \mreg/_02105_ ;
wire \mreg/_02106_ ;
wire \mreg/_02107_ ;
wire \mreg/_02108_ ;
wire \mreg/_02109_ ;
wire \mreg/_02110_ ;
wire \mreg/_02111_ ;
wire \mreg/_02112_ ;
wire \mreg/_02113_ ;
wire \mreg/_02114_ ;
wire \mreg/_02115_ ;
wire \mreg/_02116_ ;
wire \mreg/_02117_ ;
wire \mreg/_02118_ ;
wire \mreg/_02119_ ;
wire \mreg/_02120_ ;
wire \mreg/_02121_ ;
wire \mreg/_02122_ ;
wire \mreg/_02123_ ;
wire \mreg/_02124_ ;
wire \mreg/_02125_ ;
wire \mreg/_02126_ ;
wire \mreg/_02127_ ;
wire \mreg/_02128_ ;
wire \mreg/_02129_ ;
wire \mreg/_02130_ ;
wire \mreg/_02131_ ;
wire \mreg/_02132_ ;
wire \mreg/_02133_ ;
wire \mreg/_02134_ ;
wire \mreg/_02135_ ;
wire \mreg/_02136_ ;
wire \mreg/_02137_ ;
wire \mreg/_02138_ ;
wire \mreg/_02139_ ;
wire \mreg/_02140_ ;
wire \mreg/_02141_ ;
wire \mreg/_02142_ ;
wire \mreg/_02143_ ;
wire \mreg/_02144_ ;
wire \mreg/_02145_ ;
wire \mreg/_02146_ ;
wire \mreg/_02147_ ;
wire \mreg/_02148_ ;
wire \mreg/_02149_ ;
wire \mreg/_02150_ ;
wire \mreg/_02151_ ;
wire \mreg/_02152_ ;
wire \mreg/_02153_ ;
wire \mreg/_02154_ ;
wire \mreg/_02155_ ;
wire \mreg/_02156_ ;
wire \mreg/_02157_ ;
wire \mreg/_02158_ ;
wire \mreg/_02159_ ;
wire \mreg/_02160_ ;
wire \mreg/_02161_ ;
wire \mreg/_02162_ ;
wire \mreg/_02163_ ;
wire \mreg/_02164_ ;
wire \mreg/_02165_ ;
wire \mreg/_02166_ ;
wire \mreg/_02167_ ;
wire \mreg/_02168_ ;
wire \mreg/_02169_ ;
wire \mreg/_02170_ ;
wire \mreg/_02171_ ;
wire \mreg/_02172_ ;
wire \mreg/_02173_ ;
wire \mreg/_02174_ ;
wire \mreg/_02175_ ;
wire \mreg/_02176_ ;
wire \mreg/_02177_ ;
wire \mreg/_02178_ ;
wire \mreg/_02179_ ;
wire \mreg/_02180_ ;
wire \mreg/_02181_ ;
wire \mreg/_02182_ ;
wire \mreg/_02183_ ;
wire \mreg/_02184_ ;
wire \mreg/_02185_ ;
wire \mreg/_02186_ ;
wire \mreg/_02187_ ;
wire \mreg/_02188_ ;
wire \mreg/_02189_ ;
wire \mreg/_02190_ ;
wire \mreg/_02191_ ;
wire \mreg/_02192_ ;
wire \mreg/_02193_ ;
wire \mreg/_02194_ ;
wire \mreg/_02195_ ;
wire \mreg/_02196_ ;
wire \mreg/_02197_ ;
wire \mreg/_02198_ ;
wire \mreg/_02199_ ;
wire \mreg/_02200_ ;
wire \mreg/_02201_ ;
wire \mreg/_02202_ ;
wire \mreg/_02203_ ;
wire \mreg/_02204_ ;
wire \mreg/_02205_ ;
wire \mreg/_02206_ ;
wire \mreg/_02207_ ;
wire \mreg/_02208_ ;
wire \mreg/_02209_ ;
wire \mreg/_02210_ ;
wire \mreg/_02211_ ;
wire \mreg/_02212_ ;
wire \mreg/_02213_ ;
wire \mreg/_02214_ ;
wire \mreg/_02215_ ;
wire \mreg/_02216_ ;
wire \mreg/_02217_ ;
wire \mreg/_02218_ ;
wire \mreg/_02219_ ;
wire \mreg/_02220_ ;
wire \mreg/_02221_ ;
wire \mreg/_02222_ ;
wire \mreg/_02223_ ;
wire \mreg/_02224_ ;
wire \mreg/_02225_ ;
wire \mreg/_02226_ ;
wire \mreg/_02227_ ;
wire \mreg/_02228_ ;
wire \mreg/_02229_ ;
wire \mreg/_02230_ ;
wire \mreg/_02231_ ;
wire \mreg/_02232_ ;
wire \mreg/_02233_ ;
wire \mreg/_02234_ ;
wire \mreg/_02235_ ;
wire \mreg/_02236_ ;
wire \mreg/_02237_ ;
wire \mreg/_02238_ ;
wire \mreg/_02239_ ;
wire \mreg/_02240_ ;
wire \mreg/_02241_ ;
wire \mreg/_02242_ ;
wire \mreg/_02243_ ;
wire \mreg/_02244_ ;
wire \mreg/_02245_ ;
wire \mreg/_02246_ ;
wire \mreg/_02247_ ;
wire \mreg/_02248_ ;
wire \mreg/_02249_ ;
wire \mreg/_02250_ ;
wire \mreg/_02251_ ;
wire \mreg/_02252_ ;
wire \mreg/_02253_ ;
wire \mreg/_02254_ ;
wire \mreg/_02255_ ;
wire \mreg/_02256_ ;
wire \mreg/_02257_ ;
wire \mreg/_02258_ ;
wire \mreg/_02259_ ;
wire \mreg/_02260_ ;
wire \mreg/_02261_ ;
wire \mreg/_02262_ ;
wire \mreg/_02263_ ;
wire \mreg/_02264_ ;
wire \mreg/_02265_ ;
wire \mreg/_02266_ ;
wire \mreg/_02267_ ;
wire \mreg/_02268_ ;
wire \mreg/_02269_ ;
wire \mreg/_02270_ ;
wire \mreg/_02271_ ;
wire \mreg/_02272_ ;
wire \mreg/_02273_ ;
wire \mreg/_02274_ ;
wire \mreg/_02275_ ;
wire \mreg/_02276_ ;
wire \mreg/_02277_ ;
wire \mreg/_02278_ ;
wire \mreg/_02279_ ;
wire \mreg/_02280_ ;
wire \mreg/_02281_ ;
wire \mreg/_02282_ ;
wire \mreg/_02283_ ;
wire \mreg/_02284_ ;
wire \mreg/_02285_ ;
wire \mreg/_02286_ ;
wire \mreg/_02287_ ;
wire \mreg/_02288_ ;
wire \mreg/_02289_ ;
wire \mreg/_02290_ ;
wire \mreg/_02291_ ;
wire \mreg/_02292_ ;
wire \mreg/_02293_ ;
wire \mreg/_02294_ ;
wire \mreg/_02295_ ;
wire \mreg/_02296_ ;
wire \mreg/_02297_ ;
wire \mreg/_02298_ ;
wire \mreg/_02299_ ;
wire \mreg/_02300_ ;
wire \mreg/_02301_ ;
wire \mreg/_02302_ ;
wire \mreg/_02303_ ;
wire \mreg/_02304_ ;
wire \mreg/_02305_ ;
wire \mreg/_02306_ ;
wire \mreg/_02307_ ;
wire \mreg/_02308_ ;
wire \mreg/_02309_ ;
wire \mreg/_02310_ ;
wire \mreg/_02311_ ;
wire \mreg/_02312_ ;
wire \mreg/_02313_ ;
wire \mreg/_02314_ ;
wire \mreg/_02315_ ;
wire \mreg/_02316_ ;
wire \mreg/_02317_ ;
wire \mreg/_02318_ ;
wire \mreg/_02319_ ;
wire \mreg/_02320_ ;
wire \mreg/_02321_ ;
wire \mreg/_02322_ ;
wire \mreg/_02323_ ;
wire \mreg/_02324_ ;
wire \mreg/_02325_ ;
wire \mreg/_02326_ ;
wire \mreg/_02327_ ;
wire \mreg/_02328_ ;
wire \mreg/_02329_ ;
wire \mreg/_02330_ ;
wire \mreg/_02331_ ;
wire \mreg/_02332_ ;
wire \mreg/_02333_ ;
wire \mreg/_02334_ ;
wire \mreg/_02335_ ;
wire \mreg/_02336_ ;
wire \mreg/_02337_ ;
wire \mreg/_02338_ ;
wire \mreg/_02339_ ;
wire \mreg/_02340_ ;
wire \mreg/_02341_ ;
wire \mreg/_02342_ ;
wire \mreg/_02343_ ;
wire \mreg/_02344_ ;
wire \mreg/_02345_ ;
wire \mreg/_02346_ ;
wire \mreg/_02347_ ;
wire \mreg/_02348_ ;
wire \mreg/_02349_ ;
wire \mreg/_02350_ ;
wire \mreg/_02351_ ;
wire \mreg/_02352_ ;
wire \mreg/_02353_ ;
wire \mreg/_02354_ ;
wire \mreg/_02355_ ;
wire \mreg/_02356_ ;
wire \mreg/_02357_ ;
wire \mreg/_02358_ ;
wire \mreg/_02359_ ;
wire \mreg/_02360_ ;
wire \mreg/_02361_ ;
wire \mreg/_02362_ ;
wire \mreg/_02363_ ;
wire \mreg/_02364_ ;
wire \mreg/_02365_ ;
wire \mreg/_02366_ ;
wire \mreg/_02367_ ;
wire \mreg/_02368_ ;
wire \mreg/_02369_ ;
wire \mreg/_02370_ ;
wire \mreg/_02371_ ;
wire \mreg/_02372_ ;
wire \mreg/_02373_ ;
wire \mreg/_02374_ ;
wire \mreg/_02375_ ;
wire \mreg/_02376_ ;
wire \mreg/_02377_ ;
wire \mreg/_02378_ ;
wire \mreg/_02379_ ;
wire \mreg/_02380_ ;
wire \mreg/_02381_ ;
wire \mreg/_02382_ ;
wire \mreg/_02383_ ;
wire \mreg/_02384_ ;
wire \mreg/_02385_ ;
wire \mreg/_02386_ ;
wire \mreg/_02387_ ;
wire \mreg/_02388_ ;
wire \mreg/_02389_ ;
wire \mreg/_02390_ ;
wire \mreg/_02391_ ;
wire \mreg/_02392_ ;
wire \mreg/_02393_ ;
wire \mreg/_02394_ ;
wire \mreg/_02395_ ;
wire \mreg/_02396_ ;
wire \mreg/_02397_ ;
wire \mreg/_02398_ ;
wire \mreg/_02399_ ;
wire \mreg/_02400_ ;
wire \mreg/_02401_ ;
wire \mreg/_02402_ ;
wire \mreg/_02403_ ;
wire \mreg/_02404_ ;
wire \mreg/_02405_ ;
wire \mreg/_02406_ ;
wire \mreg/_02407_ ;
wire \mreg/_02408_ ;
wire \mreg/_02409_ ;
wire \mreg/_02410_ ;
wire \mreg/_02411_ ;
wire \mreg/_02412_ ;
wire \mreg/_02413_ ;
wire \mreg/_02414_ ;
wire \mreg/_02415_ ;
wire \mreg/_02416_ ;
wire \mreg/_02417_ ;
wire \mreg/_02418_ ;
wire \mreg/_02419_ ;
wire \mreg/_02420_ ;
wire \mreg/_02421_ ;
wire \mreg/_02422_ ;
wire \mreg/_02423_ ;
wire \mreg/_02424_ ;
wire \mreg/_02425_ ;
wire \mreg/_02426_ ;
wire \mreg/_02427_ ;
wire \mreg/_02428_ ;
wire \mreg/_02429_ ;
wire \mreg/_02430_ ;
wire \mreg/_02431_ ;
wire \mreg/_02432_ ;
wire \mreg/_02433_ ;
wire \mreg/_02434_ ;
wire \mreg/_02435_ ;
wire \mreg/_02436_ ;
wire \mreg/_02437_ ;
wire \mreg/_02438_ ;
wire \mreg/_02439_ ;
wire \mreg/_02440_ ;
wire \mreg/_02441_ ;
wire \mreg/_02442_ ;
wire \mreg/_02443_ ;
wire \mreg/_02444_ ;
wire \mreg/_02445_ ;
wire \mreg/_02446_ ;
wire \mreg/_02447_ ;
wire \mreg/_02448_ ;
wire \mreg/_02449_ ;
wire \mreg/_02450_ ;
wire \mreg/_02451_ ;
wire \mreg/_02452_ ;
wire \mreg/_02453_ ;
wire \mreg/_02454_ ;
wire \mreg/_02455_ ;
wire \mreg/_02456_ ;
wire \mreg/_02457_ ;
wire \mreg/_02458_ ;
wire \mreg/_02459_ ;
wire \mreg/_02460_ ;
wire \mreg/_02461_ ;
wire \mreg/_02462_ ;
wire \mreg/_02463_ ;
wire \mreg/_02464_ ;
wire \mreg/_02465_ ;
wire \mreg/_02466_ ;
wire \mreg/_02467_ ;
wire \mreg/_02468_ ;
wire \mreg/_02469_ ;
wire \mreg/_02470_ ;
wire \mreg/_02471_ ;
wire \mreg/_02472_ ;
wire \mreg/_02473_ ;
wire \mreg/_02474_ ;
wire \mreg/_02475_ ;
wire \mreg/_02476_ ;
wire \mreg/_02477_ ;
wire \mreg/_02478_ ;
wire \mreg/_02479_ ;
wire \mreg/_02480_ ;
wire \mreg/_02481_ ;
wire \mreg/_02482_ ;
wire \mreg/_02483_ ;
wire \mreg/_02484_ ;
wire \mreg/_02485_ ;
wire \mreg/_02486_ ;
wire \mreg/_02487_ ;
wire \mreg/_02488_ ;
wire \mreg/_02489_ ;
wire \mreg/_02490_ ;
wire \mreg/_02491_ ;
wire \mreg/_02492_ ;
wire \mreg/_02493_ ;
wire \mreg/_02494_ ;
wire \mreg/_02495_ ;
wire \mreg/_02496_ ;
wire \mreg/_02497_ ;
wire \mreg/_02498_ ;
wire \mreg/_02499_ ;
wire \mreg/_02500_ ;
wire \mreg/_02501_ ;
wire \mreg/_02502_ ;
wire \mreg/_02503_ ;
wire \mreg/_02504_ ;
wire \mreg/_02505_ ;
wire \mreg/_02506_ ;
wire \mreg/_02507_ ;
wire \mreg/_02508_ ;
wire \mreg/_02509_ ;
wire \mreg/_02510_ ;
wire \mreg/_02511_ ;
wire \mreg/_02512_ ;
wire \mreg/_02513_ ;
wire \mreg/_02514_ ;
wire \mreg/_02515_ ;
wire \mreg/_02516_ ;
wire \mreg/_02517_ ;
wire \mreg/_02518_ ;
wire \mreg/_02519_ ;
wire \mreg/_02520_ ;
wire \mreg/_02521_ ;
wire \mreg/_02522_ ;
wire \mreg/_02523_ ;
wire \mreg/_02524_ ;
wire \mreg/_02525_ ;
wire \mreg/_02526_ ;
wire \mreg/_02527_ ;
wire \mreg/_02528_ ;
wire \mreg/_02529_ ;
wire \mreg/_02530_ ;
wire \mreg/_02531_ ;
wire \mreg/_02532_ ;
wire \mreg/_02533_ ;
wire \mreg/_02534_ ;
wire \mreg/_02535_ ;
wire \mreg/_02536_ ;
wire \mreg/_02537_ ;
wire \mreg/_02538_ ;
wire \mreg/_02539_ ;
wire \mreg/_02540_ ;
wire \mreg/_02541_ ;
wire \mreg/_02542_ ;
wire \mreg/_02543_ ;
wire \mreg/_02544_ ;
wire \mreg/_02545_ ;
wire \mreg/_02546_ ;
wire \mreg/_02547_ ;
wire \mreg/_02548_ ;
wire \mreg/_02549_ ;
wire \mreg/_02550_ ;
wire \mreg/_02551_ ;
wire \mreg/_02552_ ;
wire \mreg/_02553_ ;
wire \mreg/_02554_ ;
wire \mreg/_02555_ ;
wire \mreg/_02556_ ;
wire \mreg/_02557_ ;
wire \mreg/_02558_ ;
wire \mreg/_02559_ ;
wire \mreg/_02560_ ;
wire \mreg/_02561_ ;
wire \mreg/_02562_ ;
wire \mreg/_02563_ ;
wire \mreg/_02564_ ;
wire \mreg/_02565_ ;
wire \mreg/_02566_ ;
wire \mreg/_02567_ ;
wire \mreg/_02568_ ;
wire \mreg/_02569_ ;
wire \mreg/_02570_ ;
wire \mreg/_02571_ ;
wire \mreg/_02572_ ;
wire \mreg/_02573_ ;
wire \mreg/_02574_ ;
wire \mreg/_02575_ ;
wire \mreg/_02576_ ;
wire \mreg/_02577_ ;
wire \mreg/_02578_ ;
wire \mreg/_02579_ ;
wire \mreg/_02580_ ;
wire \mreg/_02581_ ;
wire \mreg/_02582_ ;
wire \mreg/_02583_ ;
wire \mreg/_02584_ ;
wire \mreg/_02585_ ;
wire \mreg/_02586_ ;
wire \mreg/_02587_ ;
wire \mreg/_02588_ ;
wire \mreg/_02589_ ;
wire \mreg/_02590_ ;
wire \mreg/_02591_ ;
wire \mreg/_02592_ ;
wire \mreg/_02593_ ;
wire \mreg/_02594_ ;
wire \mreg/_02595_ ;
wire \mreg/_02596_ ;
wire \mreg/_02597_ ;
wire \mreg/_02598_ ;
wire \mreg/_02599_ ;
wire \mreg/_02600_ ;
wire \mreg/_02601_ ;
wire \mreg/_02602_ ;
wire \mreg/_02603_ ;
wire \mreg/_02604_ ;
wire \mreg/_02605_ ;
wire \mreg/_02606_ ;
wire \mreg/_02607_ ;
wire \mreg/_02608_ ;
wire \mreg/_02609_ ;
wire \mreg/_02610_ ;
wire \mreg/_02611_ ;
wire \mreg/_02612_ ;
wire \mreg/_02613_ ;
wire \mreg/_02614_ ;
wire \mreg/_02615_ ;
wire \mreg/_02616_ ;
wire \mreg/_02617_ ;
wire \mreg/_02618_ ;
wire \mreg/_02619_ ;
wire \mreg/_02620_ ;
wire \mreg/_02621_ ;
wire \mreg/_02622_ ;
wire \mreg/_02623_ ;
wire \mreg/_02624_ ;
wire \mreg/_02625_ ;
wire \mreg/_02626_ ;
wire \mreg/_02627_ ;
wire \mreg/_02628_ ;
wire \mreg/_02629_ ;
wire \mreg/_02630_ ;
wire \mreg/_02631_ ;
wire \mreg/_02632_ ;
wire \mreg/_02633_ ;
wire \mreg/_02634_ ;
wire \mreg/_02635_ ;
wire \mreg/_02636_ ;
wire \mreg/_02637_ ;
wire \mreg/_02638_ ;
wire \mreg/_02639_ ;
wire \mreg/_02640_ ;
wire \mreg/_02641_ ;
wire \mreg/_02642_ ;
wire \mreg/_02643_ ;
wire \mreg/_02644_ ;
wire \mreg/_02645_ ;
wire \mreg/_02646_ ;
wire \mreg/_02647_ ;
wire \mreg/_02648_ ;
wire \mreg/_02649_ ;
wire \mreg/_02650_ ;
wire \mreg/_02651_ ;
wire \mreg/_02652_ ;
wire \mreg/_02653_ ;
wire \mreg/_02654_ ;
wire \mreg/_02655_ ;
wire \mreg/_02656_ ;
wire \mreg/_02657_ ;
wire \mreg/_02658_ ;
wire \mreg/_02659_ ;
wire \mreg/_02660_ ;
wire \mreg/_02661_ ;
wire \mreg/_02662_ ;
wire \mreg/_02663_ ;
wire \mreg/_02664_ ;
wire \mreg/_02665_ ;
wire \mreg/_02666_ ;
wire \mreg/_02667_ ;
wire \mreg/_02668_ ;
wire \mreg/_02669_ ;
wire \mreg/_02670_ ;
wire \mreg/_02671_ ;
wire \mreg/_02672_ ;
wire \mreg/_02673_ ;
wire \mreg/_02674_ ;
wire \mreg/_02675_ ;
wire \mreg/_02676_ ;
wire \mreg/_02677_ ;
wire \mreg/_02678_ ;
wire \mreg/_02679_ ;
wire \mreg/_02680_ ;
wire \mreg/_02681_ ;
wire \mreg/_02682_ ;
wire \mreg/_02683_ ;
wire \mreg/_02684_ ;
wire \mreg/_02685_ ;
wire \mreg/_02686_ ;
wire \mreg/_02687_ ;
wire \mreg/_02688_ ;
wire \mreg/_02689_ ;
wire \mreg/_02690_ ;
wire \mreg/_02691_ ;
wire \mreg/_02692_ ;
wire \mreg/_02693_ ;
wire \mreg/_02694_ ;
wire \mreg/_02695_ ;
wire \mreg/_02696_ ;
wire \mreg/_02697_ ;
wire \mreg/_02698_ ;
wire \mreg/_02699_ ;
wire \mreg/_02700_ ;
wire \mreg/_02701_ ;
wire \mreg/_02702_ ;
wire \mreg/_02703_ ;
wire \mreg/_02704_ ;
wire \mreg/_02705_ ;
wire \mreg/_02706_ ;
wire \mreg/_02707_ ;
wire \mreg/_02708_ ;
wire \mreg/_02709_ ;
wire \mreg/_02710_ ;
wire \mreg/_02711_ ;
wire \mreg/_02712_ ;
wire \mreg/_02713_ ;
wire \mreg/_02714_ ;
wire \mreg/_02715_ ;
wire \mreg/_02716_ ;
wire \mreg/_02717_ ;
wire \mreg/_02718_ ;
wire \mreg/_02719_ ;
wire \mreg/_02720_ ;
wire \mreg/_02721_ ;
wire \mreg/_02722_ ;
wire \mreg/_02723_ ;
wire \mreg/_02724_ ;
wire \mreg/_02725_ ;
wire \mreg/_02726_ ;
wire \mreg/_02727_ ;
wire \mreg/_02728_ ;
wire \mreg/_02729_ ;
wire \mreg/_02730_ ;
wire \mreg/_02731_ ;
wire \mreg/_02732_ ;
wire \mreg/_02733_ ;
wire \mreg/_02734_ ;
wire \mreg/_02735_ ;
wire \mreg/_02736_ ;
wire \mreg/_02737_ ;
wire \mreg/_02738_ ;
wire \mreg/_02739_ ;
wire \mreg/_02740_ ;
wire \mreg/_02741_ ;
wire \mreg/_02742_ ;
wire \mreg/_02743_ ;
wire \mreg/_02744_ ;
wire \mreg/_02745_ ;
wire \mreg/_02746_ ;
wire \mreg/_02747_ ;
wire \mreg/_02748_ ;
wire \mreg/_02749_ ;
wire \mreg/_02750_ ;
wire \mreg/_02751_ ;
wire \mreg/_02752_ ;
wire \mreg/_02753_ ;
wire \mreg/_02754_ ;
wire \mreg/_02755_ ;
wire \mreg/_02756_ ;
wire \mreg/_02757_ ;
wire \mreg/_02758_ ;
wire \mreg/_02759_ ;
wire \mreg/_02760_ ;
wire \mreg/_02761_ ;
wire \mreg/_02762_ ;
wire \mreg/_02763_ ;
wire \mreg/_02764_ ;
wire \mreg/_02765_ ;
wire \mreg/_02766_ ;
wire \mreg/_02767_ ;
wire \mreg/_02768_ ;
wire \mreg/_02769_ ;
wire \mreg/_02770_ ;
wire \mreg/_02771_ ;
wire \mreg/_02772_ ;
wire \mreg/_02773_ ;
wire \mreg/_02774_ ;
wire \mreg/_02775_ ;
wire \mreg/_02776_ ;
wire \mreg/_02777_ ;
wire \mreg/_02778_ ;
wire \mreg/_02779_ ;
wire \mreg/_02780_ ;
wire \mreg/_02781_ ;
wire \mreg/_02782_ ;
wire \mreg/_02783_ ;
wire \mreg/_02784_ ;
wire \mreg/_02785_ ;
wire \mreg/_02786_ ;
wire \mreg/_02787_ ;
wire \mreg/_02788_ ;
wire \mreg/_02789_ ;
wire \mreg/_02790_ ;
wire \mreg/_02791_ ;
wire \mreg/_02792_ ;
wire \mreg/_02793_ ;
wire \mreg/_02794_ ;
wire \mreg/_02795_ ;
wire \mreg/_02796_ ;
wire \mreg/_02797_ ;
wire \mreg/_02798_ ;
wire \mreg/_02799_ ;
wire \mreg/_02800_ ;
wire \mreg/_02801_ ;
wire \mreg/_02802_ ;
wire \mreg/_02803_ ;
wire \mreg/_02804_ ;
wire \mreg/_02805_ ;
wire \mreg/_02806_ ;
wire \mreg/_02807_ ;
wire \mreg/_02808_ ;
wire \mreg/_02809_ ;
wire \mreg/_02810_ ;
wire \mreg/_02811_ ;
wire \mreg/_02812_ ;
wire \mreg/_02813_ ;
wire \mreg/_02814_ ;
wire \mreg/_02815_ ;
wire \mreg/_02816_ ;
wire \mreg/_02817_ ;
wire \mreg/_02818_ ;
wire \mreg/_02819_ ;
wire \mreg/_02820_ ;
wire \mreg/_02821_ ;
wire \mreg/_02822_ ;
wire \mreg/_02823_ ;
wire \mreg/_02824_ ;
wire \mreg/_02825_ ;
wire \mreg/_02826_ ;
wire \mreg/_02827_ ;
wire \mreg/_02828_ ;
wire \mreg/_02829_ ;
wire \mreg/_02830_ ;
wire \mreg/_02831_ ;
wire \mreg/_02832_ ;
wire \mreg/_02833_ ;
wire \mreg/_02834_ ;
wire \mreg/_02835_ ;
wire \mreg/_02836_ ;
wire \mreg/_02837_ ;
wire \mreg/_02838_ ;
wire \mreg/_02839_ ;
wire \mreg/_02840_ ;
wire \mreg/_02841_ ;
wire \mreg/_02842_ ;
wire \mreg/_02843_ ;
wire \mreg/_02844_ ;
wire \mreg/_02845_ ;
wire \mreg/_02846_ ;
wire \mreg/_02847_ ;
wire \mreg/_02848_ ;
wire \mreg/_02849_ ;
wire \mreg/_02850_ ;
wire \mreg/_02851_ ;
wire \mreg/_02852_ ;
wire \mreg/_02853_ ;
wire \mreg/_02854_ ;
wire \mreg/_02855_ ;
wire \mreg/_02856_ ;
wire \mreg/_02857_ ;
wire \mreg/_02858_ ;
wire \mreg/_02859_ ;
wire \mreg/_02860_ ;
wire \mreg/_02861_ ;
wire \mreg/_02862_ ;
wire \mreg/_02863_ ;
wire \mreg/_02864_ ;
wire \mreg/_02865_ ;
wire \mreg/_02866_ ;
wire \mreg/_02867_ ;
wire \mreg/_02868_ ;
wire \mreg/_02869_ ;
wire \mreg/_02870_ ;
wire \mreg/_02871_ ;
wire \mreg/_02872_ ;
wire \mreg/_02873_ ;
wire \mreg/_02874_ ;
wire \mreg/_02875_ ;
wire \mreg/_02876_ ;
wire \mreg/_02877_ ;
wire \mreg/_02878_ ;
wire \mreg/_02879_ ;
wire \mreg/_02880_ ;
wire \mreg/_02881_ ;
wire \mreg/_02882_ ;
wire \mreg/_02883_ ;
wire \mreg/_02884_ ;
wire \mreg/_02885_ ;
wire \mreg/_02886_ ;
wire \mreg/_02887_ ;
wire \mreg/_02888_ ;
wire \mreg/_02889_ ;
wire \mreg/_02890_ ;
wire \mreg/_02891_ ;
wire \mreg/_02892_ ;
wire \mreg/_02893_ ;
wire \mreg/_02894_ ;
wire \mreg/_02895_ ;
wire \mreg/_02896_ ;
wire \mreg/_02897_ ;
wire \mreg/_02898_ ;
wire \mreg/_02899_ ;
wire \mreg/_02900_ ;
wire \mreg/_02901_ ;
wire \mreg/_02902_ ;
wire \mreg/_02903_ ;
wire \mreg/_02904_ ;
wire \mreg/_02905_ ;
wire \mreg/_02906_ ;
wire \mreg/_02907_ ;
wire \mreg/_02908_ ;
wire \mreg/_02909_ ;
wire \mreg/_02910_ ;
wire \mreg/_02911_ ;
wire \mreg/_02912_ ;
wire \mreg/_02913_ ;
wire \mreg/_02914_ ;
wire \mreg/_02915_ ;
wire \mreg/_02916_ ;
wire \mreg/_02917_ ;
wire \mreg/_02918_ ;
wire \mreg/_02919_ ;
wire \mreg/_02920_ ;
wire \mreg/_02921_ ;
wire \mreg/_02922_ ;
wire \mreg/_02923_ ;
wire \mreg/_02924_ ;
wire \mreg/_02925_ ;
wire \mreg/_02926_ ;
wire \mreg/_02927_ ;
wire \mreg/_02928_ ;
wire \mreg/_02929_ ;
wire \mreg/_02930_ ;
wire \mreg/_02931_ ;
wire \mreg/_02932_ ;
wire \mreg/_02933_ ;
wire \mreg/_02934_ ;
wire \mreg/_02935_ ;
wire \mreg/_02936_ ;
wire \mreg/_02937_ ;
wire \mreg/_02938_ ;
wire \mreg/_02939_ ;
wire \mreg/_02940_ ;
wire \mreg/_02941_ ;
wire \mreg/_02942_ ;
wire \mreg/_02943_ ;
wire \mreg/_02944_ ;
wire \mreg/_02945_ ;
wire \mreg/_02946_ ;
wire \mreg/_02947_ ;
wire \mreg/_02948_ ;
wire \mreg/_02949_ ;
wire \mreg/_02950_ ;
wire \mreg/_02951_ ;
wire \mreg/_02952_ ;
wire \mreg/_02953_ ;
wire \mreg/_02954_ ;
wire \mreg/_02955_ ;
wire \mreg/_02956_ ;
wire \mreg/_02957_ ;
wire \mreg/_02958_ ;
wire \mreg/_02959_ ;
wire \mreg/_02960_ ;
wire \mreg/_02961_ ;
wire \mreg/_02962_ ;
wire \mreg/_02963_ ;
wire \mreg/_02964_ ;
wire \mreg/_02965_ ;
wire \mreg/_02966_ ;
wire \mreg/_02967_ ;
wire \mreg/_02968_ ;
wire \mreg/_02969_ ;
wire \mreg/_02970_ ;
wire \mreg/_02971_ ;
wire \mreg/_02972_ ;
wire \mreg/_02973_ ;
wire \mreg/_02974_ ;
wire \mreg/_02975_ ;
wire \mreg/_02976_ ;
wire \mreg/_02977_ ;
wire \mreg/_02978_ ;
wire \mreg/_02979_ ;
wire \mreg/_02980_ ;
wire \mreg/_02981_ ;
wire \mreg/_02982_ ;
wire \mreg/_02983_ ;
wire \mreg/_02984_ ;
wire \mreg/_02985_ ;
wire \mreg/_02986_ ;
wire \mreg/_02987_ ;
wire \mreg/_02988_ ;
wire \mreg/_02989_ ;
wire \mreg/_02990_ ;
wire \mreg/_02991_ ;
wire \mreg/_02992_ ;
wire \mreg/_02993_ ;
wire \mreg/_02994_ ;
wire \mreg/_02995_ ;
wire \mreg/_02996_ ;
wire \mreg/_02997_ ;
wire \mreg/_02998_ ;
wire \mreg/_02999_ ;
wire \mreg/_03000_ ;
wire \mreg/_03001_ ;
wire \mreg/_03002_ ;
wire \mreg/_03003_ ;
wire \mreg/_03004_ ;
wire \mreg/_03005_ ;
wire \mreg/_03006_ ;
wire \mreg/_03007_ ;
wire \mreg/_03008_ ;
wire \mreg/_03009_ ;
wire \mreg/_03010_ ;
wire \mreg/_03011_ ;
wire \mreg/_03012_ ;
wire \mreg/_03013_ ;
wire \mreg/_03014_ ;
wire \mreg/_03015_ ;
wire \mreg/_03016_ ;
wire \mreg/_03017_ ;
wire \mreg/_03018_ ;
wire \mreg/_03019_ ;
wire \mreg/_03020_ ;
wire \mreg/_03021_ ;
wire \mreg/_03022_ ;
wire \mreg/_03023_ ;
wire \mreg/_03024_ ;
wire \mreg/_03025_ ;
wire \mreg/_03026_ ;
wire \mreg/_03027_ ;
wire \mreg/_03028_ ;
wire \mreg/_03029_ ;
wire \mreg/_03030_ ;
wire \mreg/_03031_ ;
wire \mreg/_03032_ ;
wire \mreg/_03033_ ;
wire \mreg/_03034_ ;
wire \mreg/_03035_ ;
wire \mreg/_03036_ ;
wire \mreg/_03037_ ;
wire \mreg/_03038_ ;
wire \mreg/_03039_ ;
wire \mreg/_03040_ ;
wire \mreg/_03041_ ;
wire \mreg/_03042_ ;
wire \mreg/_03043_ ;
wire \mreg/_03044_ ;
wire \mreg/_03045_ ;
wire \mreg/_03046_ ;
wire \mreg/_03047_ ;
wire \mreg/_03048_ ;
wire \mreg/_03049_ ;
wire \mreg/_03050_ ;
wire \mreg/_03051_ ;
wire \mreg/_03052_ ;
wire \mreg/_03053_ ;
wire \mreg/_03054_ ;
wire \mreg/_03055_ ;
wire \mreg/_03056_ ;
wire \mreg/_03057_ ;
wire \mreg/_03058_ ;
wire \mreg/_03059_ ;
wire \mreg/_03060_ ;
wire \mreg/_03061_ ;
wire \mreg/_03062_ ;
wire \mreg/_03063_ ;
wire \mreg/_03064_ ;
wire \mreg/_03065_ ;
wire \mreg/_03066_ ;
wire \mreg/_03067_ ;
wire \mreg/_03068_ ;
wire \mreg/_03069_ ;
wire \mreg/_03070_ ;
wire \mreg/_03071_ ;
wire \mreg/_03072_ ;
wire \mreg/_03073_ ;
wire \mreg/_03074_ ;
wire \mreg/_03075_ ;
wire \mreg/_03076_ ;
wire \mreg/_03077_ ;
wire \mreg/_03078_ ;
wire \mreg/_03079_ ;
wire \mreg/_03080_ ;
wire \mreg/_03081_ ;
wire \mreg/_03082_ ;
wire \mreg/_03083_ ;
wire \mreg/_03084_ ;
wire \mreg/_03085_ ;
wire \mreg/_03086_ ;
wire \mreg/_03087_ ;
wire \mreg/_03088_ ;
wire \mreg/_03089_ ;
wire \mreg/_03090_ ;
wire \mreg/_03091_ ;
wire \mreg/_03092_ ;
wire \mreg/_03093_ ;
wire \mreg/_03094_ ;
wire \mreg/_03095_ ;
wire \mreg/_03096_ ;
wire \mreg/_03097_ ;
wire \mreg/_03098_ ;
wire \mreg/_03099_ ;
wire \mreg/_03100_ ;
wire \mreg/_03101_ ;
wire \mreg/_03102_ ;
wire \mreg/_03103_ ;
wire \mreg/_03104_ ;
wire \mreg/_03105_ ;
wire \mreg/_03106_ ;
wire \mreg/_03107_ ;
wire \mreg/_03108_ ;
wire \mreg/_03109_ ;
wire \mreg/_03110_ ;
wire \mreg/_03111_ ;
wire \mreg/_03112_ ;
wire \mreg/_03113_ ;
wire \mreg/_03114_ ;
wire \mreg/_03115_ ;
wire \mreg/_03116_ ;
wire \mreg/_03117_ ;
wire \mreg/_03118_ ;
wire \mreg/_03119_ ;
wire \mreg/_03120_ ;
wire \mreg/_03121_ ;
wire \mreg/_03122_ ;
wire \mreg/_03123_ ;
wire \mreg/_03124_ ;
wire \mreg/_03125_ ;
wire \mreg/_03126_ ;
wire \mreg/_03127_ ;
wire \mreg/_03128_ ;
wire \mreg/_03129_ ;
wire \mreg/_03130_ ;
wire \mreg/_03131_ ;
wire \mreg/_03132_ ;
wire \mreg/_03133_ ;
wire \mreg/_03134_ ;
wire \mreg/_03135_ ;
wire \mreg/_03136_ ;
wire \mreg/_03137_ ;
wire \mreg/_03138_ ;
wire \mreg/_03139_ ;
wire \mreg/_03140_ ;
wire \mreg/_03141_ ;
wire \mreg/_03142_ ;
wire \mreg/_03143_ ;
wire \mreg/_03144_ ;
wire \mreg/_03145_ ;
wire \mreg/_03146_ ;
wire \mreg/_03147_ ;
wire \mreg/_03148_ ;
wire \mreg/_03149_ ;
wire \mreg/_03150_ ;
wire \mreg/_03151_ ;
wire \mreg/_03152_ ;
wire \mreg/_03153_ ;
wire \mreg/_03154_ ;
wire \mreg/_03155_ ;
wire \mreg/_03156_ ;
wire \mreg/_03157_ ;
wire \mreg/_03158_ ;
wire \mreg/_03159_ ;
wire \mreg/_03160_ ;
wire \mreg/_03161_ ;
wire \mreg/_03162_ ;
wire \mreg/_03163_ ;
wire \mreg/_03164_ ;
wire \mreg/_03165_ ;
wire \mreg/_03166_ ;
wire \mreg/_03167_ ;
wire \mreg/_03168_ ;
wire \mreg/_03169_ ;
wire \mreg/_03170_ ;
wire \mreg/_03171_ ;
wire \mreg/_03172_ ;
wire \mreg/_03173_ ;
wire \mreg/_03174_ ;
wire \mreg/_03175_ ;
wire \mreg/_03176_ ;
wire \mreg/_03177_ ;
wire \mreg/_03178_ ;
wire \mreg/_03179_ ;
wire \mreg/_03180_ ;
wire \mreg/_03181_ ;
wire \mreg/_03182_ ;
wire \mreg/_03183_ ;
wire \mreg/_03184_ ;
wire \mreg/_03185_ ;
wire \mreg/_03186_ ;
wire \mreg/_03187_ ;
wire \mreg/_03188_ ;
wire \mreg/_03189_ ;
wire \mreg/_03190_ ;
wire \mreg/_03191_ ;
wire \mreg/_03192_ ;
wire \mreg/_03193_ ;
wire \mreg/_03194_ ;
wire \mreg/_03195_ ;
wire \mreg/_03196_ ;
wire \mreg/_03197_ ;
wire \mreg/_03198_ ;
wire \mreg/_03199_ ;
wire \mreg/_03200_ ;
wire \mreg/_03201_ ;
wire \mreg/_03202_ ;
wire \mreg/_03203_ ;
wire \mreg/_03204_ ;
wire \mreg/_03205_ ;
wire \mreg/_03206_ ;
wire \mreg/_03207_ ;
wire \mreg/_03208_ ;
wire \mreg/_03209_ ;
wire \mreg/_03210_ ;
wire \mreg/_03211_ ;
wire \mreg/_03212_ ;
wire \mreg/_03213_ ;
wire \mreg/_03214_ ;
wire \mreg/_03215_ ;
wire \mreg/_03216_ ;
wire \mreg/_03217_ ;
wire \mreg/_03218_ ;
wire \mreg/_03219_ ;
wire \mreg/_03220_ ;
wire \mreg/_03221_ ;
wire \mreg/_03222_ ;
wire \mreg/_03223_ ;
wire \mreg/_03224_ ;
wire \mreg/_03225_ ;
wire \mreg/_03226_ ;
wire \mreg/_03227_ ;
wire \mreg/_03228_ ;
wire \mreg/_03229_ ;
wire \mreg/_03230_ ;
wire \mreg/_03231_ ;
wire \mreg/_03232_ ;
wire \mreg/_03233_ ;
wire \mreg/_03234_ ;
wire \mreg/_03235_ ;
wire \mreg/_03236_ ;
wire \mreg/_03237_ ;
wire \mreg/_03238_ ;
wire \mreg/_03239_ ;
wire \mreg/_03240_ ;
wire \mreg/_03241_ ;
wire \mreg/_03242_ ;
wire \mreg/_03243_ ;
wire \mreg/_03244_ ;
wire \mreg/_03245_ ;
wire \mreg/_03246_ ;
wire \mreg/_03247_ ;
wire \mreg/_03248_ ;
wire \mreg/_03249_ ;
wire \mreg/_03250_ ;
wire \mreg/_03251_ ;
wire \mreg/_03252_ ;
wire \mreg/_03253_ ;
wire \mreg/_03254_ ;
wire \mreg/_03255_ ;
wire \mreg/_03256_ ;
wire \mreg/_03257_ ;
wire \mreg/_03258_ ;
wire \mreg/_03259_ ;
wire \mreg/_03260_ ;
wire \mreg/_03261_ ;
wire \mreg/_03262_ ;
wire \mreg/_03263_ ;
wire \mreg/_03264_ ;
wire \mreg/_03265_ ;
wire \mreg/_03266_ ;
wire \mreg/_03267_ ;
wire \mreg/_03268_ ;
wire \mreg/_03269_ ;
wire \mreg/_03270_ ;
wire \mreg/_03271_ ;
wire \mreg/_03272_ ;
wire \mreg/_03273_ ;
wire \mreg/_03274_ ;
wire \mreg/_03275_ ;
wire \mreg/_03276_ ;
wire \mreg/_03277_ ;
wire \mreg/_03278_ ;
wire \mreg/_03279_ ;
wire \mreg/_03280_ ;
wire \mreg/_03281_ ;
wire \mreg/_03282_ ;
wire \mreg/_03283_ ;
wire \mreg/_03284_ ;
wire \mreg/_03285_ ;
wire \mreg/_03286_ ;
wire \mreg/_03287_ ;
wire \mreg/_03288_ ;
wire \mreg/_03289_ ;
wire \mreg/_03290_ ;
wire \mreg/_03291_ ;
wire \mreg/_03292_ ;
wire \mreg/_03293_ ;
wire \mreg/_03294_ ;
wire \mreg/_03295_ ;
wire \mreg/_03296_ ;
wire \mreg/_03297_ ;
wire \mreg/_03298_ ;
wire \mreg/_03299_ ;
wire \mreg/_03300_ ;
wire \mreg/_03301_ ;
wire \mreg/_03302_ ;
wire \mreg/_03303_ ;
wire \mreg/_03304_ ;
wire \mreg/_03305_ ;
wire \mreg/_03306_ ;
wire \mreg/_03307_ ;
wire \mreg/_03308_ ;
wire \mreg/_03309_ ;
wire \mreg/_03310_ ;
wire \mreg/_03311_ ;
wire \mreg/_03312_ ;
wire \mreg/_03313_ ;
wire \mreg/_03314_ ;
wire \mreg/_03315_ ;
wire \mreg/_03316_ ;
wire \mreg/_03317_ ;
wire \mreg/_03318_ ;
wire \mreg/_03319_ ;
wire \mreg/_03320_ ;
wire \mreg/_03321_ ;
wire \mreg/_03322_ ;
wire \mreg/_03323_ ;
wire \mreg/_03324_ ;
wire \mreg/_03325_ ;
wire \mreg/_03326_ ;
wire \mreg/_03327_ ;
wire \mreg/_03328_ ;
wire \mreg/_03329_ ;
wire \mreg/_03330_ ;
wire \mreg/_03331_ ;
wire \mreg/_03332_ ;
wire \mreg/_03333_ ;
wire \mreg/_03334_ ;
wire \mreg/_03335_ ;
wire \mreg/_03336_ ;
wire \mreg/_03337_ ;
wire \mreg/_03338_ ;
wire \mreg/_03339_ ;
wire \mreg/_03340_ ;
wire \mreg/_03341_ ;
wire \mreg/_03342_ ;
wire \mreg/_03343_ ;
wire \mreg/_03344_ ;
wire \mreg/_03345_ ;
wire \mreg/_03346_ ;
wire \mreg/_03347_ ;
wire \mreg/_03348_ ;
wire \mreg/_03349_ ;
wire \mreg/_03350_ ;
wire \mreg/_03351_ ;
wire \mreg/_03352_ ;
wire \mreg/_03353_ ;
wire \mreg/_03354_ ;
wire \mreg/_03355_ ;
wire \mreg/_03356_ ;
wire \mreg/_03357_ ;
wire \mreg/_03358_ ;
wire \mreg/_03359_ ;
wire \mreg/_03360_ ;
wire \mreg/_03361_ ;
wire \mreg/_03362_ ;
wire \mreg/_03363_ ;
wire \mreg/_03364_ ;
wire \mreg/_03365_ ;
wire \mreg/_03366_ ;
wire \mreg/_03367_ ;
wire \mreg/_03368_ ;
wire \mreg/_03369_ ;
wire \mreg/_03370_ ;
wire \mreg/_03371_ ;
wire \mreg/_03372_ ;
wire \mreg/_03373_ ;
wire \mreg/_03374_ ;
wire \mreg/_03375_ ;
wire \mreg/_03376_ ;
wire \mreg/_03377_ ;
wire \mreg/_03378_ ;
wire \mreg/_03379_ ;
wire \mreg/_03380_ ;
wire \mreg/_03381_ ;
wire \mreg/_03382_ ;
wire \mreg/_03383_ ;
wire \mreg/_03384_ ;
wire \mreg/_03385_ ;
wire \mreg/_03386_ ;
wire \mreg/_03387_ ;
wire \mreg/_03388_ ;
wire \mreg/_03389_ ;
wire \mreg/_03390_ ;
wire \mreg/_03391_ ;
wire \mreg/_03392_ ;
wire \mreg/_03393_ ;
wire \mreg/_03394_ ;
wire \mreg/_03395_ ;
wire \mreg/_03396_ ;
wire \mreg/_03397_ ;
wire \mreg/_03398_ ;
wire \mreg/_03399_ ;
wire \mreg/_03400_ ;
wire \mreg/_03401_ ;
wire \mreg/_03402_ ;
wire \mreg/_03403_ ;
wire \mreg/_03404_ ;
wire \mreg/_03405_ ;
wire \mreg/_03406_ ;
wire \mreg/_03407_ ;
wire \mreg/_03408_ ;
wire \mreg/_03409_ ;
wire \mreg/_03410_ ;
wire \mreg/_03411_ ;
wire \mreg/_03412_ ;
wire \mreg/_03413_ ;
wire \mreg/_03414_ ;
wire \mreg/_03415_ ;
wire \mreg/_03416_ ;
wire \mreg/_03417_ ;
wire \mreg/_03418_ ;
wire \mreg/_03419_ ;
wire \mreg/_03420_ ;
wire \mreg/_03421_ ;
wire \mreg/_03422_ ;
wire \mreg/_03423_ ;
wire \mreg/_03424_ ;
wire \mreg/_03425_ ;
wire \mreg/_03426_ ;
wire \mreg/_03427_ ;
wire \mreg/_03428_ ;
wire \mreg/_03429_ ;
wire \mreg/_03430_ ;
wire \mreg/_03431_ ;
wire \mreg/_03432_ ;
wire \mreg/_03433_ ;
wire \mreg/_03434_ ;
wire \mreg/_03435_ ;
wire \mreg/_03436_ ;
wire \mreg/_03437_ ;
wire \mreg/_03438_ ;
wire \mreg/_03439_ ;
wire \mreg/_03440_ ;
wire \mreg/_03441_ ;
wire \mreg/_03442_ ;
wire \mreg/_03443_ ;
wire \mreg/_03444_ ;
wire \mreg/_03445_ ;
wire \mreg/_03446_ ;
wire \mreg/_03447_ ;
wire \mreg/_03448_ ;
wire \mreg/_03449_ ;
wire \mreg/_03450_ ;
wire \mreg/_03451_ ;
wire \mreg/_03452_ ;
wire \mreg/_03453_ ;
wire \mreg/_03454_ ;
wire \mreg/_03455_ ;
wire \mreg/_03456_ ;
wire \mreg/_03457_ ;
wire \mreg/_03458_ ;
wire \mreg/_03459_ ;
wire \mreg/_03460_ ;
wire \mreg/_03461_ ;
wire \mreg/_03462_ ;
wire \mreg/_03463_ ;
wire \mreg/_03464_ ;
wire \mreg/_03465_ ;
wire \mreg/_03466_ ;
wire \mreg/_03467_ ;
wire \mreg/_03468_ ;
wire \mreg/_03469_ ;
wire \mreg/_03470_ ;
wire \mreg/_03471_ ;
wire \mreg/_03472_ ;
wire \mreg/_03473_ ;
wire \mreg/_03474_ ;
wire \mreg/_03475_ ;
wire \mreg/_03476_ ;
wire \mreg/_03477_ ;
wire \mreg/_03478_ ;
wire \mreg/_03479_ ;
wire \mreg/_03480_ ;
wire \mreg/_03481_ ;
wire \mreg/_03482_ ;
wire \mreg/_03483_ ;
wire \mreg/_03484_ ;
wire \mreg/_03485_ ;
wire \mreg/_03486_ ;
wire \mreg/_03487_ ;
wire \mreg/_03488_ ;
wire \mreg/_03489_ ;
wire \mreg/_03490_ ;
wire \mreg/_03491_ ;
wire \mreg/_03492_ ;
wire \mreg/_03493_ ;
wire \mreg/_03494_ ;
wire \mreg/_03495_ ;
wire \mreg/_03496_ ;
wire \mreg/_03497_ ;
wire \mreg/_03498_ ;
wire \mreg/_03499_ ;
wire \mreg/_03500_ ;
wire \mreg/_03501_ ;
wire \mreg/_03502_ ;
wire \mreg/_03503_ ;
wire \mreg/_03504_ ;
wire \mreg/_03505_ ;
wire \mreg/_03506_ ;
wire \mreg/_03507_ ;
wire \mreg/_03508_ ;
wire \mreg/_03509_ ;
wire \mreg/_03510_ ;
wire \mreg/_03511_ ;
wire \mreg/_03512_ ;
wire \mreg/_03513_ ;
wire \mreg/_03514_ ;
wire \mreg/_03515_ ;
wire \mreg/_03516_ ;
wire \mreg/_03517_ ;
wire \mreg/_03518_ ;
wire \mreg/_03519_ ;
wire \mreg/_03520_ ;
wire \mreg/_03521_ ;
wire \mreg/_03522_ ;
wire \mreg/_03523_ ;
wire \mreg/_03524_ ;
wire \mreg/_03525_ ;
wire \mreg/_03526_ ;
wire \mreg/_03527_ ;
wire \mreg/_03528_ ;
wire \mreg/_03529_ ;
wire \mreg/_03530_ ;
wire \mreg/_03531_ ;
wire \mreg/_03532_ ;
wire \mreg/_03533_ ;
wire \mreg/_03534_ ;
wire \mreg/_03535_ ;
wire \mreg/_03536_ ;
wire \mreg/_03537_ ;
wire \mreg/_03538_ ;
wire \mreg/_03539_ ;
wire \mreg/_03540_ ;
wire \mreg/_03541_ ;
wire \mreg/_03542_ ;
wire \mreg/_03543_ ;
wire \mreg/_03544_ ;
wire \mreg/_03545_ ;
wire \mreg/_03546_ ;
wire \mreg/_03547_ ;
wire \mreg/_03548_ ;
wire \mreg/_03549_ ;
wire \mreg/_03550_ ;
wire \mreg/_03551_ ;
wire \mreg/_03552_ ;
wire \mreg/_03553_ ;
wire \mreg/_03554_ ;
wire \mreg/_03555_ ;
wire \mreg/_03556_ ;
wire \mreg/_03557_ ;
wire \mreg/_03558_ ;
wire \mreg/_03559_ ;
wire \mreg/_03560_ ;
wire \mreg/_03561_ ;
wire \mreg/_03562_ ;
wire \mreg/_03563_ ;
wire \mreg/_03564_ ;
wire \mreg/_03565_ ;
wire \mreg/_03566_ ;
wire \mreg/_03567_ ;
wire \mreg/_03568_ ;
wire \mreg/_03569_ ;
wire \mreg/_03570_ ;
wire \mreg/_03571_ ;
wire \mreg/_03572_ ;
wire \mreg/_03573_ ;
wire \mreg/_03574_ ;
wire \mreg/_03575_ ;
wire \mreg/_03576_ ;
wire \mreg/_03577_ ;
wire \mreg/_03578_ ;
wire \mreg/_03579_ ;
wire \mreg/_03580_ ;
wire \mreg/_03581_ ;
wire \mreg/_03582_ ;
wire \mreg/_03583_ ;
wire \mreg/_03584_ ;
wire \mreg/_03585_ ;
wire \mreg/_03586_ ;
wire \mreg/_03587_ ;
wire \mreg/_03588_ ;
wire \mreg/_03589_ ;
wire \mreg/_03590_ ;
wire \mreg/_03591_ ;
wire \mreg/_03592_ ;
wire \mreg/_03593_ ;
wire \mreg/_03594_ ;
wire \mreg/_03595_ ;
wire \mreg/_03596_ ;
wire \mreg/_03597_ ;
wire \mreg/_03598_ ;
wire \mreg/_03599_ ;
wire \mreg/_03600_ ;
wire \mreg/_03601_ ;
wire \mreg/_03602_ ;
wire \mreg/_03603_ ;
wire \mreg/_03604_ ;
wire \mreg/_03605_ ;
wire \mreg/_03606_ ;
wire \mreg/_03607_ ;
wire \mreg/_03608_ ;
wire \mreg/_03609_ ;
wire \mreg/_03610_ ;
wire \mreg/_03611_ ;
wire \mreg/_03612_ ;
wire \mreg/_03613_ ;
wire \mreg/_03614_ ;
wire \mreg/_03615_ ;
wire \mreg/_03616_ ;
wire \mreg/_03617_ ;
wire \mreg/_03618_ ;
wire \mreg/_03619_ ;
wire \mreg/_03620_ ;
wire \mreg/_03621_ ;
wire \mreg/_03622_ ;
wire \mreg/_03623_ ;
wire \mreg/_03624_ ;
wire \mreg/_03625_ ;
wire \mreg/_03626_ ;
wire \mreg/_03627_ ;
wire \mreg/_03628_ ;
wire \mreg/_03629_ ;
wire \mreg/_03630_ ;
wire \mreg/_03631_ ;
wire \mreg/_03632_ ;
wire \mreg/_03633_ ;
wire \mreg/_03634_ ;
wire \mreg/_03635_ ;
wire \mreg/_03636_ ;
wire \mreg/_03637_ ;
wire \mreg/_03638_ ;
wire \mreg/_03639_ ;
wire \mreg/_03640_ ;
wire \mreg/_03641_ ;
wire \mreg/_03642_ ;
wire \mreg/_03643_ ;
wire \mreg/_03644_ ;
wire \mreg/_03645_ ;
wire \mreg/_03646_ ;
wire \mreg/_03647_ ;
wire \mreg/_03648_ ;
wire \mreg/_03649_ ;
wire \mreg/_03650_ ;
wire \mreg/_03651_ ;
wire \mreg/_03652_ ;
wire \mreg/_03653_ ;
wire \mreg/_03654_ ;
wire \mreg/_03655_ ;
wire \mreg/_03656_ ;
wire \mreg/_03657_ ;
wire \mreg/_03658_ ;
wire \mreg/_03659_ ;
wire \mreg/_03660_ ;
wire \mreg/_03661_ ;
wire \mreg/_03662_ ;
wire \mreg/_03663_ ;
wire \mreg/_03664_ ;
wire \mreg/_03665_ ;
wire \mreg/_03666_ ;
wire \mreg/_03667_ ;
wire \mreg/_03668_ ;
wire \mreg/_03669_ ;
wire \mreg/_03670_ ;
wire \mreg/_03671_ ;
wire \mreg/_03672_ ;
wire \mreg/_03673_ ;
wire \mreg/_03674_ ;
wire \mreg/_03675_ ;
wire \mreg/_03676_ ;
wire \mreg/_03677_ ;
wire \mreg/_03678_ ;
wire \mreg/_03679_ ;
wire \mreg/_03680_ ;
wire \mreg/_03681_ ;
wire \mreg/_03682_ ;
wire \mreg/_03683_ ;
wire \mreg/_03684_ ;
wire \mreg/_03685_ ;
wire \mreg/_03686_ ;
wire \mreg/_03687_ ;
wire \mreg/_03688_ ;
wire \mreg/_03689_ ;
wire \mreg/_03690_ ;
wire \mreg/_03691_ ;
wire \mreg/_03692_ ;
wire \mreg/_03693_ ;
wire \mreg/_03694_ ;
wire \mreg/_03695_ ;
wire \mreg/_03696_ ;
wire \mreg/_03697_ ;
wire \mreg/_03698_ ;
wire \mreg/_03699_ ;
wire \mreg/_03700_ ;
wire \mreg/_03701_ ;
wire \mreg/_03702_ ;
wire \mreg/_03703_ ;
wire \mreg/_03704_ ;
wire \mreg/_03705_ ;
wire \mreg/_03706_ ;
wire \mreg/_03707_ ;
wire \mreg/_03708_ ;
wire \mreg/_03709_ ;
wire \mreg/_03710_ ;
wire \mreg/_03711_ ;
wire \mreg/_03712_ ;
wire \mreg/_03713_ ;
wire \mreg/_03714_ ;
wire \mreg/_03715_ ;
wire \mreg/_03716_ ;
wire \mreg/_03717_ ;
wire \mreg/_03718_ ;
wire \mreg/_03719_ ;
wire \mreg/_03720_ ;
wire \mreg/_03721_ ;
wire \mreg/_03722_ ;
wire \mreg/_03723_ ;
wire \mreg/_03724_ ;
wire \mreg/_03725_ ;
wire \mreg/_03726_ ;
wire \mreg/_03727_ ;
wire \mreg/_03728_ ;
wire \mreg/_03729_ ;
wire \mreg/_03730_ ;
wire \mreg/_03731_ ;
wire \mreg/_03732_ ;
wire \mreg/_03733_ ;
wire \mreg/_03734_ ;
wire \mreg/_03735_ ;
wire \mreg/_03736_ ;
wire \mreg/_03737_ ;
wire \mreg/_03738_ ;
wire \mreg/_03739_ ;
wire \mreg/_03740_ ;
wire \mreg/_03741_ ;
wire \mreg/_03742_ ;
wire \mreg/_03743_ ;
wire \mreg/_03744_ ;
wire \mreg/_03745_ ;
wire \mreg/_03746_ ;
wire \mreg/_03747_ ;
wire \mreg/_03748_ ;
wire \mreg/_03749_ ;
wire \mreg/_03750_ ;
wire \mreg/_03751_ ;
wire \mreg/_03752_ ;
wire \mreg/_03753_ ;
wire \mreg/_03754_ ;
wire \mreg/_03755_ ;
wire \mreg/_03756_ ;
wire \mreg/_03757_ ;
wire \mreg/_03758_ ;
wire \mreg/_03759_ ;
wire \mreg/_03760_ ;
wire \mreg/_03761_ ;
wire \mreg/_03762_ ;
wire \mreg/_03763_ ;
wire \mreg/_03764_ ;
wire \mreg/_03765_ ;
wire \mreg/_03766_ ;
wire \mreg/_03767_ ;
wire \mreg/_03768_ ;
wire \mreg/_03769_ ;
wire \mreg/_03770_ ;
wire \mreg/_03771_ ;
wire \mreg/_03772_ ;
wire \mreg/_03773_ ;
wire \mreg/_03774_ ;
wire \mreg/_03775_ ;
wire \mreg/_03776_ ;
wire \mreg/_03777_ ;
wire \mreg/_03778_ ;
wire \mreg/_03779_ ;
wire \mreg/_03780_ ;
wire \mreg/_03781_ ;
wire \mreg/_03782_ ;
wire \mreg/_03783_ ;
wire \mreg/_03784_ ;
wire \mreg/_03785_ ;
wire \mreg/_03786_ ;
wire \mreg/_03787_ ;
wire \mreg/_03788_ ;
wire \mreg/_03789_ ;
wire \mreg/_03790_ ;
wire \mreg/_03791_ ;
wire \mreg/_03792_ ;
wire \mreg/_03793_ ;
wire \mreg/_03794_ ;
wire \mreg/_03795_ ;
wire \mreg/_03796_ ;
wire \mreg/_03797_ ;
wire \mreg/_03798_ ;
wire \mreg/_03799_ ;
wire \mreg/_03800_ ;
wire \mreg/_03801_ ;
wire \mreg/_03802_ ;
wire \mreg/_03803_ ;
wire \mreg/_03804_ ;
wire \mreg/_03805_ ;
wire \mreg/_03806_ ;
wire \mreg/_03807_ ;
wire \mreg/_03808_ ;
wire \mreg/_03809_ ;
wire \mreg/_03810_ ;
wire \mreg/_03811_ ;
wire \mreg/_03812_ ;
wire \mreg/_03813_ ;
wire \mreg/_03814_ ;
wire \mreg/_03815_ ;
wire \mreg/_03816_ ;
wire \mreg/_03817_ ;
wire \mreg/_03818_ ;
wire \mreg/_03819_ ;
wire \mreg/_03820_ ;
wire \mreg/_03821_ ;
wire \mreg/_03822_ ;
wire \mreg/_03823_ ;
wire \mreg/_03824_ ;
wire \mreg/_03825_ ;
wire \mreg/_03826_ ;
wire \mreg/_03827_ ;
wire \mreg/_03828_ ;
wire \mreg/_03829_ ;
wire \mreg/_03830_ ;
wire \mreg/_03831_ ;
wire \mreg/_03832_ ;
wire \mreg/_03833_ ;
wire \mreg/_03834_ ;
wire \mreg/_03835_ ;
wire \mreg/_03836_ ;
wire \mreg/_03837_ ;
wire \mreg/_03838_ ;
wire \mreg/_03839_ ;
wire \mreg/_03840_ ;
wire \mreg/_03841_ ;
wire \mreg/_03842_ ;
wire \mreg/_03843_ ;
wire \mreg/_03844_ ;
wire \mreg/_03845_ ;
wire \mreg/_03846_ ;
wire \mreg/_03847_ ;
wire \mreg/_03848_ ;
wire \mreg/_03849_ ;
wire \mreg/_03850_ ;
wire \mreg/_03851_ ;
wire \mreg/_03852_ ;
wire \mreg/_03853_ ;
wire \mreg/_03854_ ;
wire \mreg/_03855_ ;
wire \mreg/_03856_ ;
wire \mreg/_03857_ ;
wire \mreg/_03858_ ;
wire \mreg/_03859_ ;
wire \mreg/_03860_ ;
wire \mreg/_03861_ ;
wire \mreg/_03862_ ;
wire \mreg/_03863_ ;
wire \mreg/_03864_ ;
wire \mreg/_03865_ ;
wire \mreg/_03866_ ;
wire \mreg/_03867_ ;
wire \mreg/_03868_ ;
wire \mreg/_03869_ ;
wire \mreg/_03870_ ;
wire \mreg/_03871_ ;
wire \mreg/_03872_ ;
wire \mreg/_03873_ ;
wire \mreg/_03874_ ;
wire \mreg/_03875_ ;
wire \mreg/_03876_ ;
wire \mreg/_03877_ ;
wire \mreg/_03878_ ;
wire \mreg/_03879_ ;
wire \mreg/_03880_ ;
wire \mreg/_03881_ ;
wire \mreg/_03882_ ;
wire \mreg/_03883_ ;
wire \mreg/_03884_ ;
wire \mreg/_03885_ ;
wire \mreg/_03886_ ;
wire \mreg/_03887_ ;
wire \mreg/_03888_ ;
wire \mreg/_03889_ ;
wire \mreg/_03890_ ;
wire \mreg/_03891_ ;
wire \mreg/_03892_ ;
wire \mreg/_03893_ ;
wire \mreg/_03894_ ;
wire \mreg/_03895_ ;
wire \mreg/_03896_ ;
wire \mreg/_03897_ ;
wire \mreg/_03898_ ;
wire \mreg/_03899_ ;
wire \mreg/_03900_ ;
wire \mreg/_03901_ ;
wire \mreg/_03902_ ;
wire \mreg/_03903_ ;
wire \mreg/_03904_ ;
wire \mreg/_03905_ ;
wire \mreg/_03906_ ;
wire \mreg/_03907_ ;
wire \mreg/_03908_ ;
wire \mreg/_03909_ ;
wire \mreg/_03910_ ;
wire \mreg/_03911_ ;
wire \mreg/_03912_ ;
wire \mreg/_03913_ ;
wire \mreg/_03914_ ;
wire \mreg/_03915_ ;
wire \mreg/_03916_ ;
wire \mreg/_03917_ ;
wire \mreg/_03918_ ;
wire \mreg/_03919_ ;
wire \mreg/_03920_ ;
wire \mreg/_03921_ ;
wire \mreg/_03922_ ;
wire \mreg/_03923_ ;
wire \mreg/_03924_ ;
wire \mreg/_03925_ ;
wire \mreg/_03926_ ;
wire \mreg/_03927_ ;
wire \mreg/_03928_ ;
wire \mreg/_03929_ ;
wire \mreg/_03930_ ;
wire \mreg/_03931_ ;
wire \mreg/_03932_ ;
wire \mreg/_03933_ ;
wire \mreg/_03934_ ;
wire \mreg/_03935_ ;
wire \mreg/_03936_ ;
wire \mreg/_03937_ ;
wire \mreg/_03938_ ;
wire \mreg/_03939_ ;
wire \mreg/_03940_ ;
wire \mreg/_03941_ ;
wire \mreg/_03942_ ;
wire \mreg/_03943_ ;
wire \mreg/_03944_ ;
wire \mreg/_03945_ ;
wire \mreg/_03946_ ;
wire \mreg/_03947_ ;
wire \mreg/_03948_ ;
wire \mreg/_03949_ ;
wire \mreg/_03950_ ;
wire \mreg/_03951_ ;
wire \mreg/_03952_ ;
wire \mreg/_03953_ ;
wire \mreg/_03954_ ;
wire \mreg/_03955_ ;
wire \mreg/_03956_ ;
wire \mreg/_03957_ ;
wire \mreg/_03958_ ;
wire \mreg/_03959_ ;
wire \mreg/_03960_ ;
wire \mreg/_03961_ ;
wire \mreg/_03962_ ;
wire \mreg/_03963_ ;
wire \mreg/_03964_ ;
wire \mreg/_03965_ ;
wire \mreg/_03966_ ;
wire \mreg/_03967_ ;
wire \mreg/_03968_ ;
wire \mreg/_03969_ ;
wire \mreg/_03970_ ;
wire \mreg/_03971_ ;
wire \mreg/_03972_ ;
wire \mreg/_03973_ ;
wire \mreg/_03974_ ;
wire \mreg/_03975_ ;
wire \mreg/_03976_ ;
wire \mreg/_03977_ ;
wire \mreg/_03978_ ;
wire \mreg/_03979_ ;
wire \mreg/_03980_ ;
wire \mreg/_03981_ ;
wire \mreg/_03982_ ;
wire \mreg/_03983_ ;
wire \mreg/_03984_ ;
wire \mreg/_03985_ ;
wire \mreg/_03986_ ;
wire \mreg/_03987_ ;
wire \mreg/_03988_ ;
wire \mreg/_03989_ ;
wire \mreg/_03990_ ;
wire \mreg/_03991_ ;
wire \mreg/_03992_ ;
wire \mreg/_03993_ ;
wire \mreg/_03994_ ;
wire \mreg/_03995_ ;
wire \mreg/_03996_ ;
wire \mreg/_03997_ ;
wire \mreg/_03998_ ;
wire \mreg/_03999_ ;
wire \mreg/_04000_ ;
wire \mreg/_04001_ ;
wire \mreg/_04002_ ;
wire \mreg/_04003_ ;
wire \mreg/_04004_ ;
wire \mreg/_04005_ ;
wire \mreg/_04006_ ;
wire \mreg/_04007_ ;
wire \mreg/_04008_ ;
wire \mreg/_04009_ ;
wire \mreg/_04010_ ;
wire \mreg/_04011_ ;
wire \mreg/_04012_ ;
wire \mreg/_04013_ ;
wire \mreg/_04014_ ;
wire \mreg/_04015_ ;
wire \mreg/_04016_ ;
wire \mreg/_04017_ ;
wire \mreg/_04018_ ;
wire \mreg/_04019_ ;
wire \mreg/_04020_ ;
wire \mreg/_04021_ ;
wire \mreg/_04022_ ;
wire \mreg/_04023_ ;
wire \mreg/_04024_ ;
wire \mreg/_04025_ ;
wire \mreg/_04026_ ;
wire \mreg/_04027_ ;
wire \mreg/_04028_ ;
wire \mreg/_04029_ ;
wire \mreg/_04030_ ;
wire \mreg/_04031_ ;
wire \mreg/_04032_ ;
wire \mreg/_04033_ ;
wire \mreg/_04034_ ;
wire \mreg/_04035_ ;
wire \mreg/_04036_ ;
wire \mreg/_04037_ ;
wire \mreg/_04038_ ;
wire \mreg/_04039_ ;
wire \mreg/_04040_ ;
wire \mreg/_04041_ ;
wire \mreg/_04042_ ;
wire \mreg/_04043_ ;
wire \mreg/_04044_ ;
wire \mreg/_04045_ ;
wire \mreg/_04046_ ;
wire \mreg/_04047_ ;
wire \mreg/_04048_ ;
wire \mreg/_04049_ ;
wire \mreg/_04050_ ;
wire \mreg/_04051_ ;
wire \mreg/_04052_ ;
wire \mreg/_04053_ ;
wire \mreg/_04054_ ;
wire \mreg/_04055_ ;
wire \mreg/_04056_ ;
wire \mreg/_04057_ ;
wire \mreg/_04058_ ;
wire \mreg/_04059_ ;
wire \mreg/_04060_ ;
wire \mreg/_04061_ ;
wire \mreg/_04062_ ;
wire \mreg/_04063_ ;
wire \mreg/_04064_ ;
wire \mreg/_04065_ ;
wire \mreg/_04066_ ;
wire \mreg/_04067_ ;
wire \mreg/_04068_ ;
wire \mreg/_04069_ ;
wire \mreg/_04070_ ;
wire \mreg/_04071_ ;
wire \mreg/_04072_ ;
wire \mreg/_04073_ ;
wire \mreg/_04074_ ;
wire \mreg/_04075_ ;
wire \mreg/_04076_ ;
wire \mreg/_04077_ ;
wire \mreg/_04078_ ;
wire \mreg/_04079_ ;
wire \mreg/_04080_ ;
wire \mreg/_04081_ ;
wire \mreg/_04082_ ;
wire \mreg/_04083_ ;
wire \mreg/_04084_ ;
wire \mreg/_04085_ ;
wire \mreg/_04086_ ;
wire \mreg/_04087_ ;
wire \mreg/_04088_ ;
wire \mreg/_04089_ ;
wire \mreg/_04090_ ;
wire \mreg/_04091_ ;
wire \mreg/_04092_ ;
wire \mreg/_04093_ ;
wire \mreg/_04094_ ;
wire \mreg/_04095_ ;
wire \mreg/_04096_ ;
wire \mreg/_04097_ ;
wire \mreg/_04098_ ;
wire \mreg/_04099_ ;
wire \mreg/_04100_ ;
wire \mreg/_04101_ ;
wire \mreg/_04102_ ;
wire \mreg/_04103_ ;
wire \mreg/_04104_ ;
wire \mreg/_04105_ ;
wire \mreg/_04106_ ;
wire \mreg/_04107_ ;
wire \mreg/_04108_ ;
wire \mreg/_04109_ ;
wire \mreg/_04110_ ;
wire \mreg/_04111_ ;
wire \mreg/_04112_ ;
wire \mreg/_04113_ ;
wire \mreg/_04114_ ;
wire \mreg/_04115_ ;
wire \mreg/_04116_ ;
wire \mreg/_04117_ ;
wire \mreg/_04118_ ;
wire \mreg/_04119_ ;
wire \mreg/_04120_ ;
wire \mreg/_04121_ ;
wire \mreg/_04122_ ;
wire \mreg/_04123_ ;
wire \mreg/_04124_ ;
wire \mreg/_04125_ ;
wire \mreg/_04126_ ;
wire \mreg/_04127_ ;
wire \mreg/_04128_ ;
wire \mreg/_04129_ ;
wire \mreg/_04130_ ;
wire \mreg/_04131_ ;
wire \mreg/_04132_ ;
wire \mreg/_04133_ ;
wire \mreg/_04134_ ;
wire \mreg/_04135_ ;
wire \mreg/_04136_ ;
wire \mreg/_04137_ ;
wire \mreg/_04138_ ;
wire \mreg/_04139_ ;
wire \mreg/_04140_ ;
wire \mreg/_04141_ ;
wire \mreg/_04142_ ;
wire \mreg/_04143_ ;
wire \mreg/_04144_ ;
wire \mreg/_04145_ ;
wire \mreg/_04146_ ;
wire \mreg/_04147_ ;
wire \mreg/_04148_ ;
wire \mreg/_04149_ ;
wire \mreg/_04150_ ;
wire \mreg/_04151_ ;
wire \mreg/_04152_ ;
wire \mreg/_04153_ ;
wire \mreg/_04154_ ;
wire \mreg/_04155_ ;
wire \mreg/_04156_ ;
wire \mreg/_04157_ ;
wire \mreg/_04158_ ;
wire \mreg/_04159_ ;
wire \mreg/_04160_ ;
wire \mreg/_04161_ ;
wire \mreg/_04162_ ;
wire \mreg/_04163_ ;
wire \mreg/_04164_ ;
wire \mreg/_04165_ ;
wire \mreg/_04166_ ;
wire \mreg/_04167_ ;
wire \mreg/_04168_ ;
wire \mreg/_04169_ ;
wire \mreg/_04170_ ;
wire \mreg/_04171_ ;
wire \mreg/_04172_ ;
wire \mreg/_04173_ ;
wire \mreg/_04174_ ;
wire \mreg/_04175_ ;
wire \mreg/_04176_ ;
wire \mreg/_04177_ ;
wire \mreg/_04178_ ;
wire \mreg/_04179_ ;
wire \mreg/_04180_ ;
wire \mreg/_04181_ ;
wire \mreg/_04182_ ;
wire \mreg/_04183_ ;
wire \mreg/_04184_ ;
wire \mreg/_04185_ ;
wire \mreg/_04186_ ;
wire \mreg/_04187_ ;
wire \mreg/_04188_ ;
wire \mreg/_04189_ ;
wire \mreg/_04190_ ;
wire \mreg/_04191_ ;
wire \mreg/_04192_ ;
wire \mreg/_04193_ ;
wire \mreg/_04194_ ;
wire \mreg/_04195_ ;
wire \mreg/_04196_ ;
wire \mreg/_04197_ ;
wire \mreg/_04198_ ;
wire \mreg/_04199_ ;
wire \mreg/_04200_ ;
wire \mreg/_04201_ ;
wire \mreg/_04202_ ;
wire \mreg/_04203_ ;
wire \mreg/_04204_ ;
wire \mreg/_04205_ ;
wire \mreg/_04206_ ;
wire \mreg/_04207_ ;
wire \mreg/_04208_ ;
wire \mreg/_04209_ ;
wire \mreg/_04210_ ;
wire \mreg/_04211_ ;
wire \mreg/_04212_ ;
wire \mreg/_04213_ ;
wire \mreg/_04214_ ;
wire \mreg/_04215_ ;
wire \mreg/_04216_ ;
wire \mreg/_04217_ ;
wire \mreg/_04218_ ;
wire \mreg/_04219_ ;
wire \mreg/_04220_ ;
wire \mreg/_04221_ ;
wire \mreg/_04222_ ;
wire \mreg/_04223_ ;
wire \mreg/_04224_ ;
wire \mreg/_04225_ ;
wire \mreg/_04226_ ;
wire \mreg/_04227_ ;
wire \mreg/_04228_ ;
wire \mreg/_04229_ ;
wire \mreg/_04230_ ;
wire \mreg/_04231_ ;
wire \mreg/_04232_ ;
wire \mreg/_04233_ ;
wire \mreg/_04234_ ;
wire \mreg/_04235_ ;
wire \mreg/_04236_ ;
wire \mreg/_04237_ ;
wire \mreg/_04238_ ;
wire \mreg/_04239_ ;
wire \mreg/_04240_ ;
wire \mreg/_04241_ ;
wire \mreg/_04242_ ;
wire \mreg/_04243_ ;
wire \mreg/_04244_ ;
wire \mreg/_04245_ ;
wire \mreg/_04246_ ;
wire \mreg/_04247_ ;
wire \mreg/_04248_ ;
wire \mreg/_04249_ ;
wire \mreg/_04250_ ;
wire \mreg/_04251_ ;
wire \mreg/_04252_ ;
wire \mreg/_04253_ ;
wire \mreg/_04254_ ;
wire \mreg/_04255_ ;
wire \mreg/_04256_ ;
wire \mreg/_04257_ ;
wire \mreg/_04258_ ;
wire \mreg/_04259_ ;
wire \mreg/_04260_ ;
wire \mreg/_04261_ ;
wire \mreg/_04262_ ;
wire \mreg/_04263_ ;
wire \mreg/_04264_ ;
wire \mreg/_04265_ ;
wire \mreg/_04266_ ;
wire \mreg/_04267_ ;
wire \mreg/_04268_ ;
wire \mreg/_04269_ ;
wire \mreg/_04270_ ;
wire \mreg/_04271_ ;
wire \mreg/_04272_ ;
wire \mreg/_04273_ ;
wire \mreg/_04274_ ;
wire \mreg/_04275_ ;
wire \mreg/_04276_ ;
wire \mreg/_04277_ ;
wire \mreg/_04278_ ;
wire \mreg/_04279_ ;
wire \mreg/_04280_ ;
wire \mreg/_04281_ ;
wire \mreg/_04282_ ;
wire \mreg/_04283_ ;
wire \mreg/_04284_ ;
wire \mreg/_04285_ ;
wire \mreg/_04286_ ;
wire \mreg/_04287_ ;
wire \mreg/_04288_ ;
wire \mreg/_04289_ ;
wire \mreg/_04290_ ;
wire \mreg/_04291_ ;
wire \mreg/_04292_ ;
wire \mreg/_04293_ ;
wire \mreg/_04294_ ;
wire \mreg/_04295_ ;
wire \mreg/_04296_ ;
wire \mreg/_04297_ ;
wire \mreg/_04298_ ;
wire \mreg/_04299_ ;
wire \mreg/_04300_ ;
wire \mreg/_04301_ ;
wire \mreg/_04302_ ;
wire \mreg/_04303_ ;
wire \mreg/_04304_ ;
wire \mreg/_04305_ ;
wire \mreg/_04306_ ;
wire \mreg/_04307_ ;
wire \mreg/_04308_ ;
wire \mreg/_04309_ ;
wire \mreg/_04310_ ;
wire \mreg/_04311_ ;
wire \mreg/_04312_ ;
wire \mreg/_04313_ ;
wire \mreg/_04314_ ;
wire \mreg/_04315_ ;
wire \mreg/_04316_ ;
wire \mreg/_04317_ ;
wire \mreg/_04318_ ;
wire \mreg/_04319_ ;
wire \mreg/_04320_ ;
wire \mreg/_04321_ ;
wire \mreg/_04322_ ;
wire \mreg/_04323_ ;
wire \mreg/_04324_ ;
wire \mreg/_04325_ ;
wire \mreg/_04326_ ;
wire \mreg/_04327_ ;
wire \mreg/_04328_ ;
wire \mreg/_04329_ ;
wire \mreg/_04330_ ;
wire \mreg/_04331_ ;
wire \mreg/_04332_ ;
wire \mreg/_04333_ ;
wire \mreg/_04334_ ;
wire \mreg/_04335_ ;
wire \mreg/_04336_ ;
wire \mreg/_04337_ ;
wire \mreg/_04338_ ;
wire \mreg/_04339_ ;
wire \mreg/_04340_ ;
wire \mreg/_04341_ ;
wire \mreg/_04342_ ;
wire \mreg/_04343_ ;
wire \mreg/_04344_ ;
wire \mreg/_04345_ ;
wire \mreg/_04346_ ;
wire \mreg/_04347_ ;
wire \mreg/_04348_ ;
wire \mreg/_04349_ ;
wire \mreg/_04350_ ;
wire \mreg/_04351_ ;
wire \mreg/_04352_ ;
wire \mreg/_04353_ ;
wire \mreg/_04354_ ;
wire \mreg/_04355_ ;
wire \mreg/_04356_ ;
wire \mreg/_04357_ ;
wire \mreg/_04358_ ;
wire \mreg/_04359_ ;
wire \mreg/_04360_ ;
wire \mreg/_04361_ ;
wire \mreg/_04362_ ;
wire \mreg/_04363_ ;
wire \mreg/_04364_ ;
wire \mreg/_04365_ ;
wire \mreg/_04366_ ;
wire \mreg/_04367_ ;
wire \mreg/_04368_ ;
wire \mreg/_04369_ ;
wire \mreg/_04370_ ;
wire \mreg/_04371_ ;
wire \mreg/_04372_ ;
wire \mreg/_04373_ ;
wire \mreg/_04374_ ;
wire \mreg/_04375_ ;
wire \mreg/_04376_ ;
wire \mreg/_04377_ ;
wire \mreg/_04378_ ;
wire \mreg/_04379_ ;
wire \mreg/_04380_ ;
wire \mreg/_04381_ ;
wire \mreg/_04382_ ;
wire \mreg/_04383_ ;
wire \mreg/_04384_ ;
wire \mreg/_04385_ ;
wire \mreg/_04386_ ;
wire \mreg/_04387_ ;
wire \mreg/_04388_ ;
wire \mreg/_04389_ ;
wire \mreg/_04390_ ;
wire \mreg/_04391_ ;
wire \mreg/_04392_ ;
wire \mreg/_04393_ ;
wire \mreg/_04394_ ;
wire \mreg/_04395_ ;
wire \mreg/_04396_ ;
wire \mreg/_04397_ ;
wire \mreg/_04398_ ;
wire \mreg/_04399_ ;
wire \mreg/_04400_ ;
wire \mreg/_04401_ ;
wire \mreg/_04402_ ;
wire \mreg/_04403_ ;
wire \mreg/_04404_ ;
wire \mreg/_04405_ ;
wire \mreg/_04406_ ;
wire \mreg/_04407_ ;
wire \mreg/_04408_ ;
wire \mreg/_04409_ ;
wire \mreg/_04410_ ;
wire \mreg/_04411_ ;
wire \mreg/_04412_ ;
wire \mreg/_04413_ ;
wire \mreg/_04414_ ;
wire \mreg/_04415_ ;
wire \mreg/_04416_ ;
wire \mreg/_04417_ ;
wire \mreg/_04418_ ;
wire \mreg/_04419_ ;
wire \mreg/_04420_ ;
wire \mreg/_04421_ ;
wire \mreg/_04422_ ;
wire \mreg/_04423_ ;
wire \mreg/_04424_ ;
wire \mreg/_04425_ ;
wire \mreg/_04426_ ;
wire \mreg/_04427_ ;
wire \mreg/_04428_ ;
wire \mreg/_04429_ ;
wire \mreg/_04430_ ;
wire \mreg/_04431_ ;
wire \mreg/_04432_ ;
wire \mreg/_04433_ ;
wire \mreg/_04434_ ;
wire \mreg/_04435_ ;
wire \mreg/_04436_ ;
wire \mreg/_04437_ ;
wire \mreg/_04438_ ;
wire \mreg/_04439_ ;
wire \mreg/_04440_ ;
wire \mreg/_04441_ ;
wire \mreg/_04442_ ;
wire \mreg/_04443_ ;
wire \mreg/_04444_ ;
wire \mreg/_04445_ ;
wire \mreg/_04446_ ;
wire \mreg/_04447_ ;
wire \mreg/_04448_ ;
wire \mreg/_04449_ ;
wire \mreg/_04450_ ;
wire \mreg/_04451_ ;
wire \mreg/_04452_ ;
wire \mreg/_04453_ ;
wire \mreg/_04454_ ;
wire \mreg/_04455_ ;
wire \mreg/_04456_ ;
wire \mreg/_04457_ ;
wire \mreg/_04458_ ;
wire \mreg/_04459_ ;
wire \mreg/_04460_ ;
wire \mreg/_04461_ ;
wire \mreg/_04462_ ;
wire \mreg/_04463_ ;
wire \mreg/_04464_ ;
wire \mreg/_04465_ ;
wire \mreg/_04466_ ;
wire \mreg/_04467_ ;
wire \mreg/_04468_ ;
wire \mreg/_04469_ ;
wire \mreg/_04470_ ;
wire \mreg/_04471_ ;
wire \mreg/_04472_ ;
wire \mreg/_04473_ ;
wire \mreg/_04474_ ;
wire \mreg/_04475_ ;
wire \mreg/_04476_ ;
wire \mreg/_04477_ ;
wire \mreg/_04478_ ;
wire \mreg/_04479_ ;
wire \mreg/_04480_ ;
wire \mreg/_04481_ ;
wire \mreg/_04482_ ;
wire \mreg/_04483_ ;
wire \mreg/_04484_ ;
wire \mreg/_04485_ ;
wire \mreg/_04486_ ;
wire \mreg/_04487_ ;
wire \mreg/_04488_ ;
wire \mreg/_04489_ ;
wire \mreg/_04490_ ;
wire \mreg/_04491_ ;
wire \mreg/_04492_ ;
wire \mreg/_04493_ ;
wire \mreg/_04494_ ;
wire \mreg/_04495_ ;
wire \mreg/_04496_ ;
wire \mreg/_04497_ ;
wire \mreg/_04498_ ;
wire \mreg/_04499_ ;
wire \mreg/_04500_ ;
wire \mreg/_04501_ ;
wire \mreg/_04502_ ;
wire \mreg/_04503_ ;
wire \mreg/_04504_ ;
wire \mreg/_04505_ ;
wire \mreg/_04506_ ;
wire \mreg/_04507_ ;
wire \mreg/_04508_ ;
wire \mreg/_04509_ ;
wire \mreg/_04510_ ;
wire \mreg/_04511_ ;
wire \mreg/_04512_ ;
wire \mreg/_04513_ ;
wire \mreg/_04514_ ;
wire \mreg/_04515_ ;
wire \mreg/_04516_ ;
wire \mreg/_04517_ ;
wire \mreg/_04518_ ;
wire \mreg/_04519_ ;
wire \mreg/_04520_ ;
wire \mreg/_04521_ ;
wire \mreg/_04522_ ;
wire \mreg/_04523_ ;
wire \mreg/_04524_ ;
wire \mreg/_04525_ ;
wire \mreg/_04526_ ;
wire \mreg/_04527_ ;
wire \mreg/_04528_ ;
wire \mreg/_04529_ ;
wire \mreg/_04530_ ;
wire \mreg/_04531_ ;
wire \mreg/_04532_ ;
wire \mreg/_04533_ ;
wire \mreg/_04534_ ;
wire \mreg/_04535_ ;
wire \mreg/_04536_ ;
wire \mreg/_04537_ ;
wire \mreg/_04538_ ;
wire \mreg/_04539_ ;
wire \mreg/_04540_ ;
wire \mreg/_04541_ ;
wire \mreg/_04542_ ;
wire \mreg/_04543_ ;
wire \mreg/_04544_ ;
wire \mreg/_04545_ ;
wire \mreg/_04546_ ;
wire \mreg/_04547_ ;
wire \mreg/_04548_ ;
wire \mreg/_04549_ ;
wire \mreg/_04550_ ;
wire \mreg/_04551_ ;
wire \mreg/_04552_ ;
wire \mreg/_04553_ ;
wire \mreg/_04554_ ;
wire \mreg/_04555_ ;
wire \mreg/_04556_ ;
wire \mreg/_04557_ ;
wire \mreg/_04558_ ;
wire \mreg/_04559_ ;
wire \mreg/_04560_ ;
wire \mreg/_04561_ ;
wire \mreg/_04562_ ;
wire \mreg/_04563_ ;
wire \mreg/_04564_ ;
wire \mreg/_04565_ ;
wire \mreg/_04566_ ;
wire \mreg/_04567_ ;
wire \mreg/_04568_ ;
wire \mreg/_04569_ ;
wire \mreg/_04570_ ;
wire \mreg/_04571_ ;
wire \mreg/_04572_ ;
wire \mreg/_04573_ ;
wire \mreg/_04574_ ;
wire \mreg/_04575_ ;
wire \mreg/_04576_ ;
wire \mreg/_04577_ ;
wire \mreg/_04578_ ;
wire \mreg/_04579_ ;
wire \mreg/_04580_ ;
wire \mreg/_04581_ ;
wire \mreg/_04582_ ;
wire \mreg/_04583_ ;
wire \mreg/_04584_ ;
wire \mreg/_04585_ ;
wire \mreg/_04586_ ;
wire \mreg/_04587_ ;
wire \mreg/_04588_ ;
wire \mreg/_04589_ ;
wire \mreg/_04590_ ;
wire \mreg/_04591_ ;
wire \mreg/_04592_ ;
wire \mreg/_04593_ ;
wire \mreg/_04594_ ;
wire \mreg/_04595_ ;
wire \mreg/_04596_ ;
wire \mreg/_04597_ ;
wire \mreg/_04598_ ;
wire \mreg/_04599_ ;
wire \mreg/_04600_ ;
wire \mreg/_04601_ ;
wire \mreg/_04602_ ;
wire \mreg/_04603_ ;
wire \mreg/_04604_ ;
wire \mreg/_04605_ ;
wire \mreg/_04606_ ;
wire \mreg/_04607_ ;
wire \mreg/_04608_ ;
wire \mreg/_04609_ ;
wire \mreg/_04610_ ;
wire \mreg/_04611_ ;
wire \mreg/_04612_ ;
wire \mreg/_04613_ ;
wire \mreg/_04614_ ;
wire \mreg/_04615_ ;
wire \mreg/_04616_ ;
wire \mreg/_04617_ ;
wire \mreg/_04618_ ;
wire \mreg/_04619_ ;
wire \mreg/_04620_ ;
wire \mreg/_04621_ ;
wire \mreg/_04622_ ;
wire \mreg/_04623_ ;
wire \mreg/_04624_ ;
wire \mreg/_04625_ ;
wire \mreg/_04626_ ;
wire \mreg/_04627_ ;
wire \mreg/_04628_ ;
wire \mreg/_04629_ ;
wire \mreg/_04630_ ;
wire \mreg/_04631_ ;
wire \mreg/_04632_ ;
wire \mreg/_04633_ ;
wire \mreg/_04634_ ;
wire \mreg/_04635_ ;
wire \mreg/_04636_ ;
wire \mreg/_04637_ ;
wire \mreg/_04638_ ;
wire \mreg/_04639_ ;
wire \mreg/_04640_ ;
wire \mreg/_04641_ ;
wire \mreg/_04642_ ;
wire \mreg/_04643_ ;
wire \mreg/_04644_ ;
wire \mreg/_04645_ ;
wire \mreg/_04646_ ;
wire \mreg/_04647_ ;
wire \mreg/_04648_ ;
wire \mreg/_04649_ ;
wire \mreg/_04650_ ;
wire \mreg/_04651_ ;
wire \mreg/_04652_ ;
wire \mreg/_04653_ ;
wire \mreg/_04654_ ;
wire \mreg/_04655_ ;
wire \mreg/_04656_ ;
wire \mreg/_04657_ ;
wire \mreg/_04658_ ;
wire \mreg/_04659_ ;
wire \mreg/_04660_ ;
wire \mreg/_04661_ ;
wire \mreg/_04662_ ;
wire \mreg/_04663_ ;
wire \mreg/_04664_ ;
wire \mreg/_04665_ ;
wire \mreg/_04666_ ;
wire \mreg/_04667_ ;
wire \mreg/_04668_ ;
wire \mreg/_04669_ ;
wire \mreg/_04670_ ;
wire \mreg/_04671_ ;
wire \mreg/_04672_ ;
wire \mreg/_04673_ ;
wire \mreg/_04674_ ;
wire \mreg/_04675_ ;
wire \mreg/_04676_ ;
wire \mreg/_04677_ ;
wire \mreg/_04678_ ;
wire \mreg/_04679_ ;
wire \mreg/_04680_ ;
wire \mreg/_04681_ ;
wire \mreg/_04682_ ;
wire \mreg/_04683_ ;
wire \mreg/_04684_ ;
wire \mreg/_04685_ ;
wire \mreg/_04686_ ;
wire \mreg/_04687_ ;
wire \mreg/_04688_ ;
wire \mreg/_04689_ ;
wire \mreg/_04690_ ;
wire \mreg/_04691_ ;
wire \mreg/_04692_ ;
wire \mreg/_04693_ ;
wire \mreg/_04694_ ;
wire \mreg/_04695_ ;
wire \mreg/_04696_ ;
wire \mreg/_04697_ ;
wire \mreg/_04698_ ;
wire \mreg/_04699_ ;
wire \mreg/_04700_ ;
wire \mreg/_04701_ ;
wire \mreg/_04702_ ;
wire \mreg/_04703_ ;
wire \mreg/_04704_ ;
wire \mreg/_04705_ ;
wire \mreg/_04706_ ;
wire \mreg/_04707_ ;
wire \mreg/_04708_ ;
wire \mreg/_04709_ ;
wire \mreg/_04710_ ;
wire \mreg/_04711_ ;
wire \mreg/_04712_ ;
wire \mreg/_04713_ ;
wire \mreg/_04714_ ;
wire \mreg/_04715_ ;
wire \mreg/_04716_ ;
wire \mreg/_04717_ ;
wire \mreg/_04718_ ;
wire \mreg/_04719_ ;
wire \mreg/_04720_ ;
wire \mreg/_04721_ ;
wire \mreg/_04722_ ;
wire \mreg/_04723_ ;
wire \mreg/_04724_ ;
wire \mreg/_04725_ ;
wire \mreg/_04726_ ;
wire \mreg/_04727_ ;
wire \mreg/_04728_ ;
wire \mreg/_04729_ ;
wire \mreg/_04730_ ;
wire \mreg/_04731_ ;
wire \mreg/_04732_ ;
wire \mreg/_04733_ ;
wire \mreg/_04734_ ;
wire \mreg/_04735_ ;
wire \mreg/_04736_ ;
wire \mreg/_04737_ ;
wire \mreg/_04738_ ;
wire \mreg/_04739_ ;
wire \mreg/_04740_ ;
wire \mreg/_04741_ ;
wire \mreg/_04742_ ;
wire \mreg/_04743_ ;
wire \mreg/_04744_ ;
wire \mreg/_04745_ ;
wire \mreg/_04746_ ;
wire \mreg/_04747_ ;
wire \mreg/_04748_ ;
wire \mreg/_04749_ ;
wire \mreg/_04750_ ;
wire \mreg/_04751_ ;
wire \mreg/_04752_ ;
wire \mreg/_04753_ ;
wire \mreg/_04754_ ;
wire \mreg/_04755_ ;
wire \mreg/_04756_ ;
wire \mreg/_04757_ ;
wire \mreg/_04758_ ;
wire \mreg/_04759_ ;
wire \mreg/_04760_ ;
wire \mreg/_04761_ ;
wire \mreg/_04762_ ;
wire \mreg/_04763_ ;
wire \mreg/_04764_ ;
wire \mreg/_04765_ ;
wire \mreg/_04766_ ;
wire \mreg/_04767_ ;
wire \mreg/_04768_ ;
wire \mreg/_04769_ ;
wire \mreg/_04770_ ;
wire \mreg/_04771_ ;
wire \mreg/_04772_ ;
wire \mreg/_04773_ ;
wire \mreg/_04774_ ;
wire \mreg/_04775_ ;
wire \mreg/_04776_ ;
wire \mreg/_04777_ ;
wire \mreg/_04778_ ;
wire \mreg/_04779_ ;
wire \mreg/_04780_ ;
wire \mreg/_04781_ ;
wire \mreg/_04782_ ;
wire \mreg/_04783_ ;
wire \mreg/_04784_ ;
wire \mreg/_04785_ ;
wire \mreg/_04786_ ;
wire \mreg/_04787_ ;
wire \mreg/_04788_ ;
wire \mreg/_04789_ ;
wire \mreg/_04790_ ;
wire \mreg/_04791_ ;
wire \mreg/_04792_ ;
wire \mreg/_04793_ ;
wire \mreg/_04794_ ;
wire \mreg/_04795_ ;
wire \mreg/_04796_ ;
wire \mreg/_04797_ ;
wire \mreg/_04798_ ;
wire \mreg/_04799_ ;
wire \mreg/_04800_ ;
wire \mreg/_04801_ ;
wire \mreg/_04802_ ;
wire \mreg/_04803_ ;
wire \mreg/_04804_ ;
wire \mreg/_04805_ ;
wire \mreg/_04806_ ;
wire \mreg/_04807_ ;
wire \mreg/_04808_ ;
wire \mreg/_04809_ ;
wire \mreg/_04810_ ;
wire \mreg/_04811_ ;
wire \mreg/_04812_ ;
wire \mreg/_04813_ ;
wire \mreg/_04814_ ;
wire \mreg/_04815_ ;
wire \mreg/_04816_ ;
wire \mreg/_04817_ ;
wire \mreg/_04818_ ;
wire \mreg/_04819_ ;
wire \mreg/_04820_ ;
wire \mreg/_04821_ ;
wire \mreg/_04822_ ;
wire \mreg/_04823_ ;
wire \mreg/_04824_ ;
wire \mreg/_04825_ ;
wire \mreg/_04826_ ;
wire \mreg/_04827_ ;
wire \mreg/_04828_ ;
wire \mreg/_04829_ ;
wire \mreg/_04830_ ;
wire \mreg/_04831_ ;
wire \mreg/_04832_ ;
wire \mreg/_04833_ ;
wire \mreg/_04834_ ;
wire \mreg/_04835_ ;
wire \mreg/_04836_ ;
wire \mreg/_04837_ ;
wire \mreg/_04838_ ;
wire \mreg/_04839_ ;
wire \mreg/_04840_ ;
wire \mreg/_04841_ ;
wire \mreg/_04842_ ;
wire \mreg/_04843_ ;
wire \mreg/_04844_ ;
wire \mreg/_04845_ ;
wire \mreg/_04846_ ;
wire \mreg/_04847_ ;
wire \mreg/_04848_ ;
wire \mreg/_04849_ ;
wire \mreg/_04850_ ;
wire \mreg/_04851_ ;
wire \mreg/_04852_ ;
wire \mreg/_04853_ ;
wire \mreg/_04854_ ;
wire \mreg/_04855_ ;
wire \mreg/_04856_ ;
wire \mreg/_04857_ ;
wire \mreg/_04858_ ;
wire \mreg/_04859_ ;
wire \mreg/_04860_ ;
wire \mreg/_04861_ ;
wire \mreg/_04862_ ;
wire \mreg/_04863_ ;
wire \mreg/_04864_ ;
wire \mreg/_04865_ ;
wire \mreg/_04866_ ;
wire \mreg/_04867_ ;
wire \mreg/_04868_ ;
wire \mreg/_04869_ ;
wire \mreg/_04870_ ;
wire \mreg/_04871_ ;
wire \mreg/_04872_ ;
wire \mreg/_04873_ ;
wire \mreg/_04874_ ;
wire \mreg/_04875_ ;
wire \mreg/_04876_ ;
wire \mreg/_04877_ ;
wire \mreg/_04878_ ;
wire \mreg/_04879_ ;
wire \mreg/_04880_ ;
wire \mreg/_04881_ ;
wire \mreg/_04882_ ;
wire \mreg/_04883_ ;
wire \mreg/_04884_ ;
wire \mreg/_04885_ ;
wire \mreg/_04886_ ;
wire \mreg/_04887_ ;
wire \mreg/_04888_ ;
wire \mreg/_04889_ ;
wire \mreg/_04890_ ;
wire \mreg/_04891_ ;
wire \mreg/_04892_ ;
wire \mreg/_04893_ ;
wire \mreg/_04894_ ;
wire \mreg/_04895_ ;
wire \mreg/_04896_ ;
wire \mreg/_04897_ ;
wire \mreg/_04898_ ;
wire \mreg/_04899_ ;
wire \mreg/_04900_ ;
wire \mreg/_04901_ ;
wire \mreg/_04902_ ;
wire \mreg/_04903_ ;
wire \mreg/_04904_ ;
wire \mreg/_04905_ ;
wire \mreg/_04906_ ;
wire \mreg/_04907_ ;
wire \mreg/_04908_ ;
wire \mreg/_04909_ ;
wire \mreg/_04910_ ;
wire \mreg/_04911_ ;
wire \mreg/_04912_ ;
wire \mreg/_04913_ ;
wire \mreg/_04914_ ;
wire \mreg/_04915_ ;
wire \mreg/_04916_ ;
wire \mreg/_04917_ ;
wire \mreg/_04918_ ;
wire \mreg/_04919_ ;
wire \mreg/_04920_ ;
wire \mreg/_04921_ ;
wire \mreg/_04922_ ;
wire \mreg/_04923_ ;
wire \mreg/_04924_ ;
wire \mreg/_04925_ ;
wire \mreg/_04926_ ;
wire \mreg/_04927_ ;
wire \mreg/_04928_ ;
wire \mreg/_04929_ ;
wire \mreg/_04930_ ;
wire \mreg/_04931_ ;
wire \mreg/_04932_ ;
wire \mreg/_04933_ ;
wire \mreg/_04934_ ;
wire \mreg/_04935_ ;
wire \mreg/_04936_ ;
wire \mreg/_04937_ ;
wire \mreg/_04938_ ;
wire \mreg/_04939_ ;
wire \mreg/_04940_ ;
wire \mreg/_04941_ ;
wire \mreg/_04942_ ;
wire \mreg/_04943_ ;
wire \mreg/_04944_ ;
wire \mreg/_04945_ ;
wire \mreg/_04946_ ;
wire \mreg/_04947_ ;
wire \mreg/_04948_ ;
wire \mreg/_04949_ ;
wire \mreg/_04950_ ;
wire \mreg/_04951_ ;
wire \mreg/_04952_ ;
wire \mreg/_04953_ ;
wire \mreg/_04954_ ;
wire \mreg/_04955_ ;
wire \mreg/_04956_ ;
wire \mreg/_04957_ ;
wire \mreg/_04958_ ;
wire \mreg/_04959_ ;
wire \mreg/_04960_ ;
wire \mreg/_04961_ ;
wire \mreg/_04962_ ;
wire \mreg/_04963_ ;
wire \mreg/_04964_ ;
wire \mreg/_04965_ ;
wire \mreg/_04966_ ;
wire \mreg/_04967_ ;
wire \mreg/_04968_ ;
wire \mreg/_04969_ ;
wire \mreg/_04970_ ;
wire \mreg/_04971_ ;
wire \mreg/_04972_ ;
wire \mreg/_04973_ ;
wire \mreg/_04974_ ;
wire \mreg/_04975_ ;
wire \mreg/_04976_ ;
wire \mreg/_04977_ ;
wire \mreg/_04978_ ;
wire \mreg/_04979_ ;
wire \mreg/_04980_ ;
wire \mreg/_04981_ ;
wire \mreg/_04982_ ;
wire \mreg/_04983_ ;
wire \mreg/_04984_ ;
wire \mreg/_04985_ ;
wire \mreg/_04986_ ;
wire \mreg/_04987_ ;
wire \mreg/_04988_ ;
wire \mreg/_04989_ ;
wire \mreg/_04990_ ;
wire \mreg/_04991_ ;
wire \mreg/_04992_ ;
wire \mreg/_04993_ ;
wire \mreg/_04994_ ;
wire \mreg/_04995_ ;
wire \mreg/_04996_ ;
wire \mreg/_04997_ ;
wire \mreg/_04998_ ;
wire \mreg/_04999_ ;
wire \mreg/_05000_ ;
wire \mreg/_05001_ ;
wire \mreg/_05002_ ;
wire \mreg/_05003_ ;
wire \mreg/_05004_ ;
wire \mreg/_05005_ ;
wire \mreg/_05006_ ;
wire \mreg/_05007_ ;
wire \mreg/_05008_ ;
wire \mreg/_05009_ ;
wire \mreg/_05010_ ;
wire \mreg/_05011_ ;
wire \mreg/_05012_ ;
wire \mreg/_05013_ ;
wire \mreg/_05014_ ;
wire \mreg/_05015_ ;
wire \mreg/_05016_ ;
wire \mreg/_05017_ ;
wire \mreg/_05018_ ;
wire \mreg/_05019_ ;
wire \mreg/_05020_ ;
wire \mreg/_05021_ ;
wire \mreg/_05022_ ;
wire \mreg/_05023_ ;
wire \mreg/_05024_ ;
wire \mreg/_05025_ ;
wire \mreg/_05026_ ;
wire \mreg/_05027_ ;
wire \mreg/_05028_ ;
wire \mreg/_05029_ ;
wire \mreg/_05030_ ;
wire \mreg/_05031_ ;
wire \mreg/_05032_ ;
wire \mreg/_05033_ ;
wire \mreg/_05034_ ;
wire \mreg/_05035_ ;
wire \mreg/_05036_ ;
wire \mreg/_05037_ ;
wire \mreg/_05038_ ;
wire \mreg/_05039_ ;
wire \mreg/_05040_ ;
wire \mreg/_05041_ ;
wire \mreg/_05042_ ;
wire \mreg/_05043_ ;
wire \mreg/_05044_ ;
wire \mreg/_05045_ ;
wire \mreg/_05046_ ;
wire \mreg/_05047_ ;
wire \mreg/_05048_ ;
wire \mreg/_05049_ ;
wire \mreg/_05050_ ;
wire \mreg/_05051_ ;
wire \mreg/_05052_ ;
wire \mreg/_05053_ ;
wire \mreg/_05054_ ;
wire \mreg/_05055_ ;
wire \mreg/_05056_ ;
wire \mreg/_05057_ ;
wire \mreg/_05058_ ;
wire \mreg/_05059_ ;
wire \mreg/_05060_ ;
wire \mreg/_05061_ ;
wire \mreg/_05062_ ;
wire \mreg/_05063_ ;
wire \mreg/_05064_ ;
wire \mreg/_05065_ ;
wire \mreg/_05066_ ;
wire \mreg/_05067_ ;
wire \mreg/_05068_ ;
wire \mreg/_05069_ ;
wire \mreg/_05070_ ;
wire \mreg/_05071_ ;
wire \mreg/_05072_ ;
wire \mreg/_05073_ ;
wire \mreg/_05074_ ;
wire \mreg/_05075_ ;
wire \mreg/_05076_ ;
wire \mreg/_05077_ ;
wire \mreg/_05078_ ;
wire \mreg/_05079_ ;
wire \mreg/_05080_ ;
wire \mreg/_05081_ ;
wire \mreg/_05082_ ;
wire \mreg/_05083_ ;
wire \mreg/_05084_ ;
wire \mreg/_05085_ ;
wire \mreg/_05086_ ;
wire \mreg/_05087_ ;
wire \mreg/_05088_ ;
wire \mreg/_05089_ ;
wire \mreg/_05090_ ;
wire \mreg/_05091_ ;
wire \mreg/_05092_ ;
wire \mreg/_05093_ ;
wire \mreg/_05094_ ;
wire \mreg/_05095_ ;
wire \mreg/_05096_ ;
wire \mreg/_05097_ ;
wire \mreg/_05098_ ;
wire \mreg/_05099_ ;
wire \mreg/_05100_ ;
wire \mreg/_05101_ ;
wire \mreg/_05102_ ;
wire \mreg/_05103_ ;
wire \mreg/_05104_ ;
wire \mreg/_05105_ ;
wire \mreg/_05106_ ;
wire \mreg/_05107_ ;
wire \mreg/_05108_ ;
wire \mreg/_05109_ ;
wire \mreg/_05110_ ;
wire \mreg/_05111_ ;
wire \mreg/_05112_ ;
wire \mreg/_05113_ ;
wire \mreg/_05114_ ;
wire \mreg/_05115_ ;
wire \mreg/_05116_ ;
wire \mreg/_05117_ ;
wire \mreg/_05118_ ;
wire \mreg/_05119_ ;
wire \mreg/_05120_ ;
wire \mreg/_05121_ ;
wire \mreg/_05122_ ;
wire \mreg/_05123_ ;
wire \mreg/_05124_ ;
wire \mreg/_05125_ ;
wire \mreg/_05126_ ;
wire \mreg/_05127_ ;
wire \mreg/_05128_ ;
wire \mreg/_05129_ ;
wire \mreg/_05130_ ;
wire \mreg/_05131_ ;
wire \mreg/_05132_ ;
wire \mreg/_05133_ ;
wire \mreg/_05134_ ;
wire \mreg/_05135_ ;
wire \mreg/_05136_ ;
wire \mreg/_05137_ ;
wire \mreg/_05138_ ;
wire \mreg/_05139_ ;
wire \mreg/_05140_ ;
wire \mreg/_05141_ ;
wire \mreg/_05142_ ;
wire \mreg/_05143_ ;
wire \mreg/_05144_ ;
wire \mreg/_05145_ ;
wire \mreg/_05146_ ;
wire \mreg/_05147_ ;
wire \mreg/_05148_ ;
wire \mreg/_05149_ ;
wire \mreg/_05150_ ;
wire \mreg/_05151_ ;
wire \mreg/_05152_ ;
wire \mreg/_05153_ ;
wire \mreg/_05154_ ;
wire \mreg/_05155_ ;
wire \mreg/_05156_ ;
wire \mreg/_05157_ ;
wire \mreg/_05158_ ;
wire \mreg/_05159_ ;
wire \mreg/_05160_ ;
wire \mreg/_05161_ ;
wire \mreg/_05162_ ;
wire \mreg/_05163_ ;
wire \mreg/_05164_ ;
wire \mreg/_05165_ ;
wire \mreg/_05166_ ;
wire \mreg/_05167_ ;
wire \mreg/_05168_ ;
wire \mreg/_05169_ ;
wire \mreg/_05170_ ;
wire \mreg/_05171_ ;
wire \mreg/_05172_ ;
wire \mreg/_05173_ ;
wire \mreg/_05174_ ;
wire \mreg/_05175_ ;
wire \mreg/_05176_ ;
wire \mreg/_05177_ ;
wire \mreg/_05178_ ;
wire \mreg/_05179_ ;
wire \mreg/_05180_ ;
wire \mreg/_05181_ ;
wire \mreg/_05182_ ;
wire \mreg/_05183_ ;
wire \mreg/_05184_ ;
wire \mreg/_05185_ ;
wire \mreg/_05186_ ;
wire \mreg/_05187_ ;
wire \mreg/_05188_ ;
wire \mreg/_05189_ ;
wire \mreg/_05190_ ;
wire \mreg/_05191_ ;
wire \mreg/_05192_ ;
wire \mreg/_05193_ ;
wire \mreg/_05194_ ;
wire \mreg/_05195_ ;
wire \mreg/_05196_ ;
wire \mreg/_05197_ ;
wire \mreg/_05198_ ;
wire \mreg/_05199_ ;
wire \mreg/_05200_ ;
wire \mreg/_05201_ ;
wire \mreg/_05202_ ;
wire \mreg/_05203_ ;
wire \mreg/_05204_ ;
wire \mreg/_05205_ ;
wire \mreg/_05206_ ;
wire \mreg/_05207_ ;
wire \mreg/_05208_ ;
wire \mreg/_05209_ ;
wire \mreg/_05210_ ;
wire \mreg/_05211_ ;
wire \mreg/_05212_ ;
wire \mreg/_05213_ ;
wire \mreg/_05214_ ;
wire \mreg/_05215_ ;
wire \mreg/_05216_ ;
wire \mreg/_05217_ ;
wire \mreg/_05218_ ;
wire \mreg/_05219_ ;
wire \mreg/_05220_ ;
wire \mreg/_05221_ ;
wire \mreg/_05222_ ;
wire \mreg/_05223_ ;
wire \mreg/_05224_ ;
wire \mreg/_05225_ ;
wire \mreg/_05226_ ;
wire \mreg/_05227_ ;
wire \mreg/_05228_ ;
wire \mreg/_05229_ ;
wire \mreg/_05230_ ;
wire \mreg/_05231_ ;
wire \mreg/_05232_ ;
wire \mreg/_05233_ ;
wire \mreg/_05234_ ;
wire \mreg/_05235_ ;
wire \mreg/_05236_ ;
wire \mreg/_05237_ ;
wire \mreg/_05238_ ;
wire \mreg/_05239_ ;
wire \mreg/_05240_ ;
wire \mreg/_05241_ ;
wire \mreg/_05242_ ;
wire \mreg/_05243_ ;
wire \mreg/_05244_ ;
wire \mreg/_05245_ ;
wire \mreg/_05246_ ;
wire \mreg/_05247_ ;
wire \mreg/_05248_ ;
wire \mreg/_05249_ ;
wire \mreg/_05250_ ;
wire \mreg/_05251_ ;
wire \mreg/_05252_ ;
wire \mreg/_05253_ ;
wire \mreg/_05254_ ;
wire \mreg/_05255_ ;
wire \mreg/_05256_ ;
wire \mreg/_05257_ ;
wire \mreg/_05258_ ;
wire \mreg/_05259_ ;
wire \mreg/_05260_ ;
wire \mreg/_05261_ ;
wire \mreg/_05262_ ;
wire \mreg/_05263_ ;
wire \mreg/_05264_ ;
wire \mreg/_05265_ ;
wire \mreg/_05266_ ;
wire \mreg/_05267_ ;
wire \mreg/_05268_ ;
wire \mreg/_05269_ ;
wire \mreg/_05270_ ;
wire \mreg/_05271_ ;
wire \mreg/_05272_ ;
wire \mreg/_05273_ ;
wire \mreg/_05274_ ;
wire \mreg/_05275_ ;
wire \mreg/_05276_ ;
wire \mreg/_05277_ ;
wire \mreg/_05278_ ;
wire \mreg/_05279_ ;
wire \mreg/_05280_ ;
wire \mreg/_05281_ ;
wire \mreg/_05282_ ;
wire \mreg/_05283_ ;
wire \mreg/_05284_ ;
wire \mreg/_05285_ ;
wire \mreg/_05286_ ;
wire \mreg/_05287_ ;
wire \mreg/_05288_ ;
wire \mreg/_05289_ ;
wire \mreg/_05290_ ;
wire \mreg/_05291_ ;
wire \mreg/_05292_ ;
wire \mreg/_05293_ ;
wire \mreg/_05294_ ;
wire \mreg/_05295_ ;
wire \mreg/_05296_ ;
wire \mreg/_05297_ ;
wire \mreg/_05298_ ;
wire \mreg/_05299_ ;
wire \mreg/_05300_ ;
wire \mreg/_05301_ ;
wire \mreg/_05302_ ;
wire \mreg/_05303_ ;
wire \mreg/_05304_ ;
wire \mreg/_05305_ ;
wire \mreg/_05306_ ;
wire \mreg/_05307_ ;
wire \mreg/_05308_ ;
wire \mreg/_05309_ ;
wire \mreg/_05310_ ;
wire \mreg/_05311_ ;
wire \mreg/_05312_ ;
wire \mreg/_05313_ ;
wire \mreg/_05314_ ;
wire \mreg/_05315_ ;
wire \mreg/_05316_ ;
wire \mreg/_05317_ ;
wire \mreg/_05318_ ;
wire \mreg/_05319_ ;
wire \mreg/_05320_ ;
wire \mreg/_05321_ ;
wire \mreg/_05322_ ;
wire \mreg/_05323_ ;
wire \mreg/_05324_ ;
wire \mreg/_05325_ ;
wire \mreg/_05326_ ;
wire \mreg/_05327_ ;
wire \mreg/_05328_ ;
wire \mreg/_05329_ ;
wire \mreg/_05330_ ;
wire \mreg/_05331_ ;
wire \mreg/_05332_ ;
wire \mreg/_05333_ ;
wire \mreg/_05334_ ;
wire \mreg/_05335_ ;
wire \mreg/_05336_ ;
wire \mreg/_05337_ ;
wire \mreg/_05338_ ;
wire \mreg/_05339_ ;
wire \mreg/_05340_ ;
wire \mreg/_05341_ ;
wire \mreg/_05342_ ;
wire \mreg/_05343_ ;
wire \mreg/_05344_ ;
wire \mreg/_05345_ ;
wire \mreg/_05346_ ;
wire \mreg/_05347_ ;
wire \mreg/_05348_ ;
wire \mreg/_05349_ ;
wire \mreg/_05350_ ;
wire \mreg/_05351_ ;
wire \mreg/_05352_ ;
wire \mreg/_05353_ ;
wire \mreg/_05354_ ;
wire \mreg/_05355_ ;
wire \mreg/_05356_ ;
wire \mreg/_05357_ ;
wire \mreg/_05358_ ;
wire \mreg/_05359_ ;
wire \mreg/_05360_ ;
wire \mreg/_05361_ ;
wire \mreg/_05362_ ;
wire \mreg/_05363_ ;
wire \mreg/_05364_ ;
wire \mreg/_05365_ ;
wire \mreg/_05366_ ;
wire \mreg/_05367_ ;
wire \mreg/_05368_ ;
wire \mreg/_05369_ ;
wire \mreg/_05370_ ;
wire \mreg/_05371_ ;
wire \mreg/_05372_ ;
wire \mreg/_05373_ ;
wire \mreg/_05374_ ;
wire \mreg/_05375_ ;
wire \mreg/_05376_ ;
wire \mreg/_05377_ ;
wire \mreg/_05378_ ;
wire \mreg/_05379_ ;
wire \mreg/_05380_ ;
wire \mreg/_05381_ ;
wire \mreg/_05382_ ;
wire \mreg/_05383_ ;
wire \mreg/_05384_ ;
wire \mreg/_05385_ ;
wire \mreg/_05386_ ;
wire \mreg/_05387_ ;
wire \mreg/_05388_ ;
wire \mreg/_05389_ ;
wire \mreg/_05390_ ;
wire \mreg/_05391_ ;
wire \mreg/_05392_ ;
wire \mreg/_05393_ ;
wire \mreg/_05394_ ;
wire \mreg/_05395_ ;
wire \mreg/_05396_ ;
wire \mreg/_05397_ ;
wire \mreg/_05398_ ;
wire \mreg/_05399_ ;
wire \mreg/_05400_ ;
wire \mreg/_05401_ ;
wire \mreg/_05402_ ;
wire \mreg/_05403_ ;
wire \mreg/_05404_ ;
wire \mreg/_05405_ ;
wire \mreg/_05406_ ;
wire \mreg/_05407_ ;
wire \mreg/_05408_ ;
wire \mreg/_05409_ ;
wire \mreg/_05410_ ;
wire \mreg/_05411_ ;
wire \mreg/_05412_ ;
wire \mreg/_05413_ ;
wire \mreg/_05414_ ;
wire \mreg/_05415_ ;
wire \mreg/_05416_ ;
wire \mreg/_05417_ ;
wire \mreg/_05418_ ;
wire \mreg/_05419_ ;
wire \mreg/_05420_ ;
wire \mreg/_05421_ ;
wire \mreg/_05422_ ;
wire \mreg/_05423_ ;
wire \mreg/_05424_ ;
wire \mreg/_05425_ ;
wire \mreg/_05426_ ;
wire \mreg/_05427_ ;
wire \mreg/_05428_ ;
wire \mreg/_05429_ ;
wire \mreg/_05430_ ;
wire \mreg/_05431_ ;
wire \mreg/_05432_ ;
wire \mreg/_05433_ ;
wire \mreg/_05434_ ;
wire \mreg/_05435_ ;
wire \mreg/_05436_ ;
wire \mreg/_05437_ ;
wire \mreg/_05438_ ;
wire \mreg/_05439_ ;
wire \mreg/_05440_ ;
wire \mreg/_05441_ ;
wire \mreg/_05442_ ;
wire \mreg/_05443_ ;
wire \mreg/_05444_ ;
wire \mreg/_05445_ ;
wire \mreg/_05446_ ;
wire \mreg/_05447_ ;
wire \mreg/_05448_ ;
wire \mreg/_05449_ ;
wire \mreg/_05450_ ;
wire \mreg/_05451_ ;
wire \mreg/_05452_ ;
wire \mreg/_05453_ ;
wire \mreg/_05454_ ;
wire \mreg/_05455_ ;
wire \mreg/_05456_ ;
wire \mreg/_05457_ ;
wire \mreg/_05458_ ;
wire \mreg/_05459_ ;
wire \mreg/_05460_ ;
wire \mreg/_05461_ ;
wire \mreg/_05462_ ;
wire \mreg/_05463_ ;
wire \mreg/_05464_ ;
wire \mreg/_05465_ ;
wire \mreg/_05466_ ;
wire \mreg/_05467_ ;
wire \mreg/_05468_ ;
wire \mreg/_05469_ ;
wire \mreg/_05470_ ;
wire \mreg/_05471_ ;
wire \mreg/_05472_ ;
wire \mreg/_05473_ ;
wire \mreg/_05474_ ;
wire \mreg/_05475_ ;
wire \mreg/_05476_ ;
wire \mreg/_05477_ ;
wire \mreg/_05478_ ;
wire \mreg/_05479_ ;
wire \mreg/_05480_ ;
wire \mreg/_05481_ ;
wire \mreg/_05482_ ;
wire \mreg/_05483_ ;
wire \mreg/_05484_ ;
wire \mreg/_05485_ ;
wire \mreg/_05486_ ;
wire \mreg/_05487_ ;
wire \mreg/_05488_ ;
wire \mreg/_05489_ ;
wire \mreg/_05490_ ;
wire \mreg/_05491_ ;
wire \mreg/_05492_ ;
wire \mreg/_05493_ ;
wire \mreg/_05494_ ;
wire \mreg/_05495_ ;
wire \mreg/_05496_ ;
wire \mreg/_05497_ ;
wire \mreg/_05498_ ;
wire \mreg/_05499_ ;
wire \mreg/_05500_ ;
wire \mreg/_05501_ ;
wire \mreg/_05502_ ;
wire \mreg/_05503_ ;
wire \mreg/_05504_ ;
wire \mreg/_05505_ ;
wire \mreg/_05506_ ;
wire \mreg/_05507_ ;
wire \mreg/_05508_ ;
wire \mreg/_05509_ ;
wire \mreg/_05510_ ;
wire \mreg/_05511_ ;
wire \mreg/_05512_ ;
wire \mreg/_05513_ ;
wire \mreg/_05514_ ;
wire \mreg/_05515_ ;
wire \mreg/_05516_ ;
wire \mreg/_05517_ ;
wire \mreg/_05518_ ;
wire \mreg/_05519_ ;
wire \mreg/_05520_ ;
wire \mreg/_05521_ ;
wire \mreg/_05522_ ;
wire \mreg/_05523_ ;
wire \mreg/_05524_ ;
wire \mreg/_05525_ ;
wire \mreg/_05526_ ;
wire \mreg/_05527_ ;
wire \mreg/_05528_ ;
wire \mreg/_05529_ ;
wire \mreg/_05530_ ;
wire \mreg/_05531_ ;
wire \mreg/_05532_ ;
wire \mreg/_05533_ ;
wire \mreg/_05534_ ;
wire \mreg/_05535_ ;
wire \mreg/_05536_ ;
wire \mreg/_05537_ ;
wire \mreg/_05538_ ;
wire \mreg/_05539_ ;
wire \mreg/_05540_ ;
wire \mreg/_05541_ ;
wire \mreg/_05542_ ;
wire \mreg/_05543_ ;
wire \mreg/_05544_ ;
wire \mreg/_05545_ ;
wire \mreg/_05546_ ;
wire \mreg/_05547_ ;
wire \mreg/_05548_ ;
wire \mreg/_05549_ ;
wire \mreg/_05550_ ;
wire \mreg/_05551_ ;
wire \mreg/_05552_ ;
wire \mreg/_05553_ ;
wire \mreg/_05554_ ;
wire \mreg/_05555_ ;
wire \mreg/_05556_ ;
wire \mreg/_05557_ ;
wire \mreg/_05558_ ;
wire \mreg/_05559_ ;
wire \mreg/_05560_ ;
wire \mreg/_05561_ ;
wire \mreg/_05562_ ;
wire \mreg/_05563_ ;
wire \mreg/_05564_ ;
wire \mreg/_05565_ ;
wire \mreg/_05566_ ;
wire \mreg/_05567_ ;
wire \mreg/_05568_ ;
wire \mreg/_05569_ ;
wire \mreg/_05570_ ;
wire \mreg/_05571_ ;
wire \mreg/_05572_ ;
wire \mreg/_05573_ ;
wire \mreg/_05574_ ;
wire \mreg/_05575_ ;
wire \mreg/_05576_ ;
wire \mreg/_05577_ ;
wire \mreg/_05578_ ;
wire \mreg/_05579_ ;
wire \mreg/_05580_ ;
wire \mreg/_05581_ ;
wire \mreg/_05582_ ;
wire \mreg/_05583_ ;
wire \mreg/_05584_ ;
wire \mreg/_05585_ ;
wire \mreg/_05586_ ;
wire \mreg/_05587_ ;
wire \mreg/_05588_ ;
wire \mreg/_05589_ ;
wire \mreg/_05590_ ;
wire \mreg/_05591_ ;
wire \mreg/_05592_ ;
wire \mreg/_05593_ ;
wire \mreg/_05594_ ;
wire \mreg/_05595_ ;
wire \mreg/_05596_ ;
wire \mreg/_05597_ ;
wire \mreg/_05598_ ;
wire \mreg/_05599_ ;
wire \mreg/_05600_ ;
wire \mreg/_05601_ ;
wire \mreg/_05602_ ;
wire \mreg/_05603_ ;
wire \mreg/_05604_ ;
wire \mreg/_05605_ ;
wire \mreg/_05606_ ;
wire \mreg/_05607_ ;
wire \mreg/_05608_ ;
wire \mreg/_05609_ ;
wire \mreg/_05610_ ;
wire \mreg/_05611_ ;
wire \mreg/_05612_ ;
wire \mreg/_05613_ ;
wire \mreg/_05614_ ;
wire \mreg/_05615_ ;
wire \mreg/_05616_ ;
wire \mreg/_05617_ ;
wire \mreg/_05618_ ;
wire \mreg/_05619_ ;
wire \mreg/_05620_ ;
wire \mreg/_05621_ ;
wire \mreg/_05622_ ;
wire \mreg/_05623_ ;
wire \mreg/_05624_ ;
wire \mreg/_05625_ ;
wire \mreg/_05626_ ;
wire \mreg/_05627_ ;
wire \mreg/_05628_ ;
wire \mreg/_05629_ ;
wire \mreg/_05630_ ;
wire \mreg/_05631_ ;
wire \mreg/_05632_ ;
wire \mreg/_05633_ ;
wire \mreg/_05634_ ;
wire \mreg/_05635_ ;
wire \mreg/_05636_ ;
wire \mreg/_05637_ ;
wire \mreg/_05638_ ;
wire \mreg/_05639_ ;
wire \mreg/_05640_ ;
wire \mreg/_05641_ ;
wire \mreg/_05642_ ;
wire \mreg/_05643_ ;
wire \mreg/_05644_ ;
wire \mreg/_05645_ ;
wire \mreg/_05646_ ;
wire \mreg/_05647_ ;
wire \mreg/_05648_ ;
wire \mreg/_05649_ ;
wire \mreg/_05650_ ;
wire \mreg/_05651_ ;
wire \mreg/_05652_ ;
wire \mreg/_05653_ ;
wire \mreg/_05654_ ;
wire \mreg/_05655_ ;
wire \mreg/_05656_ ;
wire \mreg/_05657_ ;
wire \mreg/_05658_ ;
wire \mreg/_05659_ ;
wire \mreg/_05660_ ;
wire \mreg/_05661_ ;
wire \mreg/_05662_ ;
wire \mreg/_05663_ ;
wire \mreg/_05664_ ;
wire \mreg/_05665_ ;
wire \mreg/_05666_ ;
wire \mreg/_05667_ ;
wire \mreg/_05668_ ;
wire \mreg/_05669_ ;
wire \mreg/_05670_ ;
wire \mreg/_05671_ ;
wire \mreg/_05672_ ;
wire \mreg/_05673_ ;
wire \mreg/_05674_ ;
wire \mreg/_05675_ ;
wire \mreg/_05676_ ;
wire \mreg/_05677_ ;
wire \mreg/_05678_ ;
wire \mreg/_05679_ ;
wire \mreg/_05680_ ;
wire \mreg/_05681_ ;
wire \mreg/_05682_ ;
wire \mreg/_05683_ ;
wire \mreg/_05684_ ;
wire \mreg/_05685_ ;
wire \mreg/_05686_ ;
wire \mreg/_05687_ ;
wire \mreg/_05688_ ;
wire \mreg/_05689_ ;
wire \mreg/_05690_ ;
wire \mreg/_05691_ ;
wire \mreg/_05692_ ;
wire \mreg/_05693_ ;
wire \mreg/_05694_ ;
wire \mreg/_05695_ ;
wire \mreg/_05696_ ;
wire \mreg/_05697_ ;
wire \mreg/_05698_ ;
wire \mreg/_05699_ ;
wire \mreg/_05700_ ;
wire \mreg/_05701_ ;
wire \mreg/_05702_ ;
wire \mreg/_05703_ ;
wire \mreg/_05704_ ;
wire \mreg/_05705_ ;
wire \mreg/_05706_ ;
wire \mreg/_05707_ ;
wire \mreg/_05708_ ;
wire \mreg/_05709_ ;
wire \mreg/_05710_ ;
wire \mreg/_05711_ ;
wire \mreg/_05712_ ;
wire \mreg/_05713_ ;
wire \mreg/_05714_ ;
wire \mreg/_05715_ ;
wire \mreg/_05716_ ;
wire \mreg/_05717_ ;
wire \mreg/_05718_ ;
wire \mreg/_05719_ ;
wire \mreg/_05720_ ;
wire \mreg/_05721_ ;
wire \mreg/_05722_ ;
wire \mreg/_05723_ ;
wire \mreg/_05724_ ;
wire \mreg/_05725_ ;
wire \mreg/_05726_ ;
wire \mreg/_05727_ ;
wire \mreg/_05728_ ;
wire \mreg/_05729_ ;
wire \mreg/_05730_ ;
wire \mreg/_05731_ ;
wire \mreg/_05732_ ;
wire \mreg/_05733_ ;
wire \mreg/_05734_ ;
wire \mreg/_05735_ ;
wire \mreg/_05736_ ;
wire \mreg/_05737_ ;
wire \mreg/_05738_ ;
wire \mreg/_05739_ ;
wire \mreg/_05740_ ;
wire \mreg/_05741_ ;
wire \mreg/_05742_ ;
wire \mreg/_05743_ ;
wire \mreg/_05744_ ;
wire \mreg/_05745_ ;
wire \mreg/_05746_ ;
wire \mreg/_05747_ ;
wire \mreg/_05748_ ;
wire \mreg/_05749_ ;
wire \mreg/_05750_ ;
wire \mreg/_05751_ ;
wire \mreg/_05752_ ;
wire \mreg/_05753_ ;
wire \mreg/_05754_ ;
wire \mreg/_05755_ ;
wire \mreg/_05756_ ;
wire \mreg/_05757_ ;
wire \mreg/_05758_ ;
wire \mreg/_05759_ ;
wire \mreg/_05760_ ;
wire \mreg/_05761_ ;
wire \mreg/_05762_ ;
wire \mreg/_05763_ ;
wire \mreg/_05764_ ;
wire \mreg/_05765_ ;
wire \mreg/_05766_ ;
wire \mreg/_05767_ ;
wire \mreg/_05768_ ;
wire \mreg/_05769_ ;
wire \mreg/_05770_ ;
wire \mreg/_05771_ ;
wire \mreg/_05772_ ;
wire \mreg/_05773_ ;
wire \mreg/_05774_ ;
wire \mreg/_05775_ ;
wire \mreg/_05776_ ;
wire \mreg/_05777_ ;
wire \mreg/_05778_ ;
wire \mreg/_05779_ ;
wire \mreg/_05780_ ;
wire \mreg/_05781_ ;
wire \mreg/_05782_ ;
wire \mreg/_05783_ ;
wire \mreg/_05784_ ;
wire \mreg/_05785_ ;
wire \mreg/_05786_ ;
wire \mreg/_05787_ ;
wire \mreg/_05788_ ;
wire \mreg/_05789_ ;
wire \mreg/_05790_ ;
wire \mreg/_05791_ ;
wire \mreg/_05792_ ;
wire \mreg/_05793_ ;
wire \mreg/_05794_ ;
wire \mreg/_05795_ ;
wire \mreg/_05796_ ;
wire \mreg/_05797_ ;
wire \mreg/_05798_ ;
wire \mreg/_05799_ ;
wire \mreg/_05800_ ;
wire \mreg/_05801_ ;
wire \mreg/_05802_ ;
wire \mreg/_05803_ ;
wire \mreg/_05804_ ;
wire \mreg/_05805_ ;
wire \mreg/_05806_ ;
wire \mreg/_05807_ ;
wire \mreg/_05808_ ;
wire \mreg/_05809_ ;
wire \mreg/_05810_ ;
wire \mreg/_05811_ ;
wire \mreg/_05812_ ;
wire \mreg/_05813_ ;
wire \mreg/_05814_ ;
wire \mreg/_05815_ ;
wire \mreg/_05816_ ;
wire \mreg/_05817_ ;
wire \mreg/_05818_ ;
wire \mreg/_05819_ ;
wire \mreg/_05820_ ;
wire \mreg/_05821_ ;
wire \mreg/_05822_ ;
wire \mreg/_05823_ ;
wire \mreg/_05824_ ;
wire \mreg/_05825_ ;
wire \mreg/_05826_ ;
wire \mreg/_05827_ ;
wire \mreg/_05828_ ;
wire \mreg/_05829_ ;
wire \mreg/_05830_ ;
wire \mreg/_05831_ ;
wire \mreg/_05832_ ;
wire \mreg/_05833_ ;
wire \mreg/_05834_ ;
wire \mreg/_05835_ ;
wire \mreg/_05836_ ;
wire \mreg/_05837_ ;
wire \mreg/_05838_ ;
wire \mreg/_05839_ ;
wire \mreg/_05840_ ;
wire \mreg/_05841_ ;
wire \mreg/_05842_ ;
wire \mreg/_05843_ ;
wire \mreg/_05844_ ;
wire \mreg/_05845_ ;
wire \mreg/_05846_ ;
wire \mreg/_05847_ ;
wire \mreg/_05848_ ;
wire \mreg/_05849_ ;
wire \mreg/_05850_ ;
wire \mreg/_05851_ ;
wire \mreg/_05852_ ;
wire \mreg/_05853_ ;
wire \mreg/_05854_ ;
wire \mreg/_05855_ ;
wire \mreg/_05856_ ;
wire \mreg/_05857_ ;
wire \mreg/_05858_ ;
wire \mreg/_05859_ ;
wire \mreg/_05860_ ;
wire \mreg/_05861_ ;
wire \mreg/_05862_ ;
wire \mreg/_05863_ ;
wire \mreg/_05864_ ;
wire \mreg/_05865_ ;
wire \mreg/_05866_ ;
wire \mreg/_05867_ ;
wire \mreg/_05868_ ;
wire \mreg/_05869_ ;
wire \mreg/_05870_ ;
wire \mreg/_05871_ ;
wire \mreg/_05872_ ;
wire \mreg/_05873_ ;
wire \mreg/_05874_ ;
wire \mreg/_05875_ ;
wire \mreg/_05876_ ;
wire \mreg/_05877_ ;
wire \mreg/_05878_ ;
wire \mreg/_05879_ ;
wire \mreg/_05880_ ;
wire \mreg/_05881_ ;
wire \mreg/_05882_ ;
wire \mreg/_05883_ ;
wire \mreg/_05884_ ;
wire \mreg/_05885_ ;
wire \mreg/_05886_ ;
wire \mreg/_05887_ ;
wire \mreg/_05888_ ;
wire \mreg/_05889_ ;
wire \mreg/_05890_ ;
wire \mreg/_05891_ ;
wire \mreg/_05892_ ;
wire \mreg/_05893_ ;
wire \mreg/_05894_ ;
wire \mreg/_05895_ ;
wire \mreg/_05896_ ;
wire \mreg/_05897_ ;
wire \mreg/_05898_ ;
wire \mreg/_05899_ ;
wire \mreg/_05900_ ;
wire \mreg/_05901_ ;
wire \mreg/_05902_ ;
wire \mreg/_05903_ ;
wire \mreg/_05904_ ;
wire \mreg/_05905_ ;
wire \mreg/_05906_ ;
wire \mreg/_05907_ ;
wire \mreg/_05908_ ;
wire \mreg/_05909_ ;
wire \mreg/_05910_ ;
wire \mreg/_05911_ ;
wire \mreg/_05912_ ;
wire \mreg/_05913_ ;
wire \mreg/_05914_ ;
wire \mreg/_05915_ ;
wire \mreg/_05916_ ;
wire \mreg/_05917_ ;
wire \mreg/_05918_ ;
wire \mreg/_05919_ ;
wire \mreg/_05920_ ;
wire \mreg/_05921_ ;
wire \mreg/_05922_ ;
wire \mreg/_05923_ ;
wire \mreg/_05924_ ;
wire \mreg/_05925_ ;
wire \mreg/_05926_ ;
wire \mreg/_05927_ ;
wire \mreg/_05928_ ;
wire \mreg/_05929_ ;
wire \mreg/_05930_ ;
wire \mreg/_05931_ ;
wire \mreg/_05932_ ;
wire \mreg/_05933_ ;
wire \mreg/_05934_ ;
wire \mreg/_05935_ ;
wire \mreg/_05936_ ;
wire \mreg/_05937_ ;
wire \mreg/_05938_ ;
wire \mreg/_05939_ ;
wire \mreg/_05940_ ;
wire \mreg/_05941_ ;
wire \mreg/_05942_ ;
wire \mreg/_05943_ ;
wire \mreg/_05944_ ;
wire \mreg/_05945_ ;
wire \mreg/_05946_ ;
wire \mreg/_05947_ ;
wire \mreg/_05948_ ;
wire \mreg/_05949_ ;
wire \mreg/_05950_ ;
wire \mreg/_05951_ ;
wire \mreg/_05952_ ;
wire \mreg/_05953_ ;
wire \mreg/_05954_ ;
wire \mreg/_05955_ ;
wire \mreg/_05956_ ;
wire \mreg/_05957_ ;
wire \mreg/_05958_ ;
wire \mreg/_05959_ ;
wire \mreg/_05960_ ;
wire \mreg/_05961_ ;
wire \mreg/_05962_ ;
wire \mreg/_05963_ ;
wire \mreg/_05964_ ;
wire \mreg/_05965_ ;
wire \mreg/_05966_ ;
wire \mreg/_05967_ ;
wire \mreg/_05968_ ;
wire \mreg/_05969_ ;
wire \mreg/_05970_ ;
wire \mreg/_05971_ ;
wire \mreg/_05972_ ;
wire \mreg/_05973_ ;
wire \mreg/_05974_ ;
wire \mreg/_05975_ ;
wire \mreg/_05976_ ;
wire \mreg/_05977_ ;
wire \mreg/_05978_ ;
wire \mreg/_05979_ ;
wire \mreg/_05980_ ;
wire \mreg/_05981_ ;
wire \mreg/_05982_ ;
wire \mreg/_05983_ ;
wire \mreg/_05984_ ;
wire \mreg/_05985_ ;
wire \mreg/_05986_ ;
wire \mreg/_05987_ ;
wire \mreg/_05988_ ;
wire \mreg/_05989_ ;
wire \mreg/_05990_ ;
wire \mreg/_05991_ ;
wire \mreg/_05992_ ;
wire \mreg/_05993_ ;
wire \mreg/_05994_ ;
wire \mreg/_05995_ ;
wire \mreg/_05996_ ;
wire \mreg/_05997_ ;
wire \mreg/_05998_ ;
wire \mreg/_05999_ ;
wire \mreg/_06000_ ;
wire \mreg/_06001_ ;
wire \mreg/_06002_ ;
wire \mreg/_06003_ ;
wire \mreg/_06004_ ;
wire \mreg/_06005_ ;
wire \mreg/_06006_ ;
wire \mreg/_06007_ ;
wire \mreg/_06008_ ;
wire \mreg/_06009_ ;
wire \mreg/_06010_ ;
wire \mreg/_06011_ ;
wire \mreg/_06012_ ;
wire \mreg/_06013_ ;
wire \mreg/_06014_ ;
wire \mreg/_06015_ ;
wire \mreg/_06016_ ;
wire \mreg/_06017_ ;
wire \mreg/_06018_ ;
wire \mreg/_06019_ ;
wire \mreg/_06020_ ;
wire \mreg/_06021_ ;
wire \mreg/_06022_ ;
wire \mreg/_06023_ ;
wire \mreg/_06024_ ;
wire \mreg/_06025_ ;
wire \mreg/_06026_ ;
wire \mreg/_06027_ ;
wire \mreg/_06028_ ;
wire \mreg/_06029_ ;
wire \mreg/_06030_ ;
wire \mreg/_06031_ ;
wire \mreg/_06032_ ;
wire \mreg/_06033_ ;
wire \mreg/_06034_ ;
wire \mreg/_06035_ ;
wire \mreg/_06036_ ;
wire \mreg/_06037_ ;
wire \mreg/_06038_ ;
wire \mreg/_06039_ ;
wire \mreg/_06040_ ;
wire \mreg/_06041_ ;
wire \mreg/_06042_ ;
wire \mreg/_06043_ ;
wire \mreg/_06044_ ;
wire \mreg/_06045_ ;
wire \mreg/_06046_ ;
wire \mreg/_06047_ ;
wire \mreg/_06048_ ;
wire \mreg/_06049_ ;
wire \mreg/_06050_ ;
wire \mreg/_06051_ ;
wire \mreg/_06052_ ;
wire \mreg/_06053_ ;
wire \mreg/_06054_ ;
wire \mreg/_06055_ ;
wire \mreg/_06056_ ;
wire \mreg/_06057_ ;
wire \mreg/_06058_ ;
wire \mreg/_06059_ ;
wire \mreg/_06060_ ;
wire \mreg/_06061_ ;
wire \mreg/_06062_ ;
wire \mreg/_06063_ ;
wire \mreg/_06064_ ;
wire \mreg/_06065_ ;
wire \mreg/_06066_ ;
wire \mreg/_06067_ ;
wire \mreg/_06068_ ;
wire \mreg/_06069_ ;
wire \mreg/_06070_ ;
wire \mreg/_06071_ ;
wire \mreg/_06072_ ;
wire \mreg/_06073_ ;
wire \mreg/_06074_ ;
wire \mreg/_06075_ ;
wire \mreg/_06076_ ;
wire \mreg/_06077_ ;
wire \mreg/_06078_ ;
wire \mreg/_06079_ ;
wire \mreg/_06080_ ;
wire \mreg/_06081_ ;
wire \mreg/_06082_ ;
wire \mreg/_06083_ ;
wire \mreg/_06084_ ;
wire \mreg/_06085_ ;
wire \mreg/_06086_ ;
wire \mreg/_06087_ ;
wire \mreg/_06088_ ;
wire \mreg/_06089_ ;
wire \mreg/_06090_ ;
wire \mreg/_06091_ ;
wire \mreg/_06092_ ;
wire \mreg/_06093_ ;
wire \mreg/_06094_ ;
wire \mreg/_06095_ ;
wire \mreg/_06096_ ;
wire \mreg/_06097_ ;
wire \mreg/_06098_ ;
wire \mreg/_06099_ ;
wire \mreg/_06100_ ;
wire \mreg/_06101_ ;
wire \mreg/_06102_ ;
wire \mreg/_06103_ ;
wire \mreg/_06104_ ;
wire \mreg/_06105_ ;
wire \mreg/_06106_ ;
wire \mreg/_06107_ ;
wire \mreg/_06108_ ;
wire \mreg/_06109_ ;
wire \mreg/_06110_ ;
wire \mreg/_06111_ ;
wire \mreg/_06112_ ;
wire \mreg/_06113_ ;
wire \mreg/_06114_ ;
wire \mreg/_06115_ ;
wire \mreg/_06116_ ;
wire \mreg/_06117_ ;
wire \mreg/_06118_ ;
wire \mreg/_06119_ ;
wire \mreg/_06120_ ;
wire \mreg/_06121_ ;
wire \mreg/_06122_ ;
wire \mreg/_06123_ ;
wire \mreg/_06124_ ;
wire \mreg/_06125_ ;
wire \mreg/_06126_ ;
wire \mreg/_06127_ ;
wire \mreg/_06128_ ;
wire \mreg/_06129_ ;
wire \mreg/_06130_ ;
wire \mreg/_06131_ ;
wire \mreg/_06132_ ;
wire \mreg/_06133_ ;
wire \mreg/_06134_ ;
wire \mreg/_06135_ ;
wire \mreg/_06136_ ;
wire \mreg/_06137_ ;
wire \mreg/_06138_ ;
wire \mreg/_06139_ ;
wire \mreg/_06140_ ;
wire \mreg/_06141_ ;
wire \mreg/_06142_ ;
wire \mreg/_06143_ ;
wire \mreg/_06144_ ;
wire \mreg/_06145_ ;
wire \mreg/_06146_ ;
wire \mreg/_06147_ ;
wire \mreg/_06148_ ;
wire \mreg/_06149_ ;
wire \mreg/_06150_ ;
wire \mreg/_06151_ ;
wire \mreg/_06152_ ;
wire \mreg/_06153_ ;
wire \mreg/_06154_ ;
wire \mreg/_06155_ ;
wire \mreg/_06156_ ;
wire \mreg/_06157_ ;
wire \mreg/_06158_ ;
wire \mreg/_06159_ ;
wire \mreg/_06160_ ;
wire \mreg/_06161_ ;
wire \mreg/_06162_ ;
wire \mreg/_06163_ ;
wire \mreg/_06164_ ;
wire \mreg/_06165_ ;
wire \mreg/_06166_ ;
wire \mreg/_06167_ ;
wire \mreg/_06168_ ;
wire \mreg/_06169_ ;
wire \mreg/_06170_ ;
wire \mreg/_06171_ ;
wire \mreg/_06172_ ;
wire \mreg/_06173_ ;
wire \mreg/_06174_ ;
wire \mreg/_06175_ ;
wire \mreg/_06176_ ;
wire \mreg/_06177_ ;
wire \mreg/_06178_ ;
wire \mreg/_06179_ ;
wire \mreg/_06180_ ;
wire \mreg/_06181_ ;
wire \mreg/_06182_ ;
wire \mreg/_06183_ ;
wire \mreg/_06184_ ;
wire \mreg/_06185_ ;
wire \mreg/_06186_ ;
wire \mreg/_06187_ ;
wire \mreg/_06188_ ;
wire \mreg/_06189_ ;
wire \mreg/_06190_ ;
wire \mreg/_06191_ ;
wire \mreg/_06192_ ;
wire \mreg/_06193_ ;
wire \mreg/_06194_ ;
wire \mreg/_06195_ ;
wire \mreg/_06196_ ;
wire \mreg/_06197_ ;
wire \mreg/_06198_ ;
wire \mreg/_06199_ ;
wire \mreg/_06200_ ;
wire \mreg/_06201_ ;
wire \mreg/_06202_ ;
wire \mreg/_06203_ ;
wire \mreg/_06204_ ;
wire \mreg/_06205_ ;
wire \mreg/_06206_ ;
wire \mreg/_06207_ ;
wire \mreg/_06208_ ;
wire \mreg/_06209_ ;
wire \mreg/_06210_ ;
wire \mreg/_06211_ ;
wire \mreg/_06212_ ;
wire \mreg/_06213_ ;
wire \mreg/_06214_ ;
wire \mreg/_06215_ ;
wire \mreg/_06216_ ;
wire \mreg/_06217_ ;
wire \mreg/_06218_ ;
wire \mreg/_06219_ ;
wire \mreg/_06220_ ;
wire \mreg/_06221_ ;
wire \mreg/_06222_ ;
wire \mreg/_06223_ ;
wire \mreg/_06224_ ;
wire \mreg/_06225_ ;
wire \mreg/_06226_ ;
wire \mreg/_06227_ ;
wire \mreg/_06228_ ;
wire \mreg/_06229_ ;
wire \mreg/_06230_ ;
wire \mreg/_06231_ ;
wire \mreg/_06232_ ;
wire \mreg/_06233_ ;
wire \mreg/_06234_ ;
wire \mreg/_06235_ ;
wire \mreg/_06236_ ;
wire \mreg/_06237_ ;
wire \mreg/_06238_ ;
wire \mreg/_06239_ ;
wire \mreg/_06240_ ;
wire \mreg/_06241_ ;
wire \mreg/_06242_ ;
wire \mreg/_06243_ ;
wire \mreg/_06244_ ;
wire \mreg/_06245_ ;
wire \mreg/_06246_ ;
wire \mreg/_06247_ ;
wire \mreg/_06248_ ;
wire \mreg/_06249_ ;
wire \mreg/_06250_ ;
wire \mreg/_06251_ ;
wire \mreg/_06252_ ;
wire \mreg/_06253_ ;
wire \mreg/_06254_ ;
wire \mreg/_06255_ ;
wire \mreg/_06256_ ;
wire \mreg/_06257_ ;
wire \mreg/_06258_ ;
wire \mreg/_06259_ ;
wire \mreg/_06260_ ;
wire \mreg/_06261_ ;
wire \mreg/_06262_ ;
wire \mreg/_06263_ ;
wire \mreg/_06264_ ;
wire \mreg/_06265_ ;
wire \mreg/_06266_ ;
wire \mreg/_06267_ ;
wire \mreg/_06268_ ;
wire \mreg/_06269_ ;
wire \mreg/_06270_ ;
wire \mreg/_06271_ ;
wire \mreg/_06272_ ;
wire \mreg/_06273_ ;
wire \mreg/_06274_ ;
wire \mreg/_06275_ ;
wire \mreg/_06276_ ;
wire \mreg/_06277_ ;
wire \mreg/_06278_ ;
wire \mreg/_06279_ ;
wire \mreg/_06280_ ;
wire \mreg/_06281_ ;
wire \mreg/_06282_ ;
wire \mreg/_06283_ ;
wire \mreg/_06284_ ;
wire \mreg/_06285_ ;
wire \mreg/_06286_ ;
wire \mreg/_06287_ ;
wire \mreg/_06288_ ;
wire \mreg/_06289_ ;
wire \mreg/_06290_ ;
wire \mreg/_06291_ ;
wire \mreg/_06292_ ;
wire \mreg/_06293_ ;
wire \mreg/_06294_ ;
wire \mreg/_06295_ ;
wire \mreg/_06296_ ;
wire \mreg/_06297_ ;
wire \mreg/_06298_ ;
wire \mreg/_06299_ ;
wire \mreg/_06300_ ;
wire \mreg/_06301_ ;
wire \mreg/_06302_ ;
wire \mreg/_06303_ ;
wire \mreg/_06304_ ;
wire \mreg/_06305_ ;
wire \mreg/_06306_ ;
wire \mreg/_06307_ ;
wire \mreg/_06308_ ;
wire \mreg/_06309_ ;
wire \mreg/_06310_ ;
wire \mreg/_06311_ ;
wire \mreg/_06312_ ;
wire \mreg/_06313_ ;
wire \mreg/_06314_ ;
wire \mreg/_06315_ ;
wire \mreg/_06316_ ;
wire \mreg/_06317_ ;
wire \mreg/_06318_ ;
wire \mreg/_06319_ ;
wire \mreg/_06320_ ;
wire \mreg/_06321_ ;
wire \mreg/_06322_ ;
wire \mreg/_06323_ ;
wire \mreg/_06324_ ;
wire \mreg/_06325_ ;
wire \mreg/_06326_ ;
wire \mreg/_06327_ ;
wire \mreg/_06328_ ;
wire \mreg/_06329_ ;
wire \mreg/_06330_ ;
wire \mreg/_06331_ ;
wire \mreg/_06332_ ;
wire \mreg/_06333_ ;
wire \mreg/_06334_ ;
wire \mreg/_06335_ ;
wire \mreg/_06336_ ;
wire \mreg/_06337_ ;
wire \mreg/_06338_ ;
wire \mreg/_06339_ ;
wire \mreg/_06340_ ;
wire \mreg/_06341_ ;
wire \mreg/_06342_ ;
wire \mreg/_06343_ ;
wire \mreg/_06344_ ;
wire \mreg/_06345_ ;
wire \mreg/_06346_ ;
wire \mreg/_06347_ ;
wire \mreg/_06348_ ;
wire \mreg/_06349_ ;
wire \mreg/_06350_ ;
wire \mreg/_06351_ ;
wire \mreg/_06352_ ;
wire \mreg/_06353_ ;
wire \mreg/_06354_ ;
wire \mreg/_06355_ ;
wire \mreg/_06356_ ;
wire \mreg/_06357_ ;
wire \mreg/_06358_ ;
wire \mreg/_06359_ ;
wire \mreg/_06360_ ;
wire \mreg/_06361_ ;
wire \mreg/_06362_ ;
wire \mreg/_06363_ ;
wire \mreg/_06364_ ;
wire \mreg/_06365_ ;
wire \mreg/_06366_ ;
wire \mreg/_06367_ ;
wire \mreg/_06368_ ;
wire \mreg/_06369_ ;
wire \mreg/_06370_ ;
wire \mreg/_06371_ ;
wire \mreg/_06372_ ;
wire \mreg/_06373_ ;
wire \mreg/_06374_ ;
wire \mreg/_06375_ ;
wire \mreg/_06376_ ;
wire \mreg/_06377_ ;
wire \mreg/_06378_ ;
wire \mreg/_06379_ ;
wire \mreg/_06380_ ;
wire \mreg/_06381_ ;
wire \mreg/_06382_ ;
wire \mreg/_06383_ ;
wire \mreg/_06384_ ;
wire \mreg/_06385_ ;
wire \mreg/_06386_ ;
wire \mreg/_06387_ ;
wire \mreg/_06388_ ;
wire \mreg/_06389_ ;
wire \mreg/_06390_ ;
wire \mreg/_06391_ ;
wire \mreg/_06392_ ;
wire \mreg/_06393_ ;
wire \mreg/_06394_ ;
wire \mreg/_06395_ ;
wire \mreg/_06396_ ;
wire \mreg/_06397_ ;
wire \mreg/_06398_ ;
wire \mreg/_06399_ ;
wire \mreg/_06400_ ;
wire \mreg/_06401_ ;
wire \mreg/_06402_ ;
wire \mreg/_06403_ ;
wire \mreg/_06404_ ;
wire \mreg/_06405_ ;
wire \mreg/_06406_ ;
wire \mreg/_06407_ ;
wire \mreg/_06408_ ;
wire \mreg/_06409_ ;
wire \mreg/_06410_ ;
wire \mreg/_06411_ ;
wire \mreg/_06412_ ;
wire \mreg/_06413_ ;
wire \mreg/_06414_ ;
wire \mreg/_06415_ ;
wire \mreg/_06416_ ;
wire \mreg/_06417_ ;
wire \mreg/_06418_ ;
wire \mreg/_06419_ ;
wire \mreg/_06420_ ;
wire \mreg/_06421_ ;
wire \mreg/_06422_ ;
wire \mreg/_06423_ ;
wire \mreg/_06424_ ;
wire \mreg/_06425_ ;
wire \mreg/_06426_ ;
wire \mreg/_06427_ ;
wire \mreg/_06428_ ;
wire \mreg/_06429_ ;
wire \mreg/_06430_ ;
wire \mreg/_06431_ ;
wire \mreg/_06432_ ;
wire \mreg/_06433_ ;
wire \mreg/_06434_ ;
wire \mreg/_06435_ ;
wire \mreg/_06436_ ;
wire \mreg/_06437_ ;
wire \mreg/_06438_ ;
wire \mreg/_06439_ ;
wire \mreg/_06440_ ;
wire \mreg/_06441_ ;
wire \mreg/_06442_ ;
wire \mreg/_06443_ ;
wire \mreg/_06444_ ;
wire \mreg/_06445_ ;
wire \mreg/_06446_ ;
wire \mreg/_06447_ ;
wire \mreg/_06448_ ;
wire \mreg/_06449_ ;
wire \mreg/_06450_ ;
wire \mreg/_06451_ ;
wire \mreg/_06452_ ;
wire \mreg/_06453_ ;
wire \mreg/_06454_ ;
wire \mreg/_06455_ ;
wire \mreg/_06456_ ;
wire \mreg/_06457_ ;
wire \mreg/_06458_ ;
wire \mreg/_06459_ ;
wire \mreg/_06460_ ;
wire \mreg/_06461_ ;
wire \mreg/_06462_ ;
wire \mreg/_06463_ ;
wire \mreg/_06464_ ;
wire \mreg/_06465_ ;
wire \mreg/_06466_ ;
wire \mreg/_06467_ ;
wire \mreg/_06468_ ;
wire \mreg/_06469_ ;
wire \mreg/_06470_ ;
wire \mreg/_06471_ ;
wire \mreg/_06472_ ;
wire \mreg/_06473_ ;
wire \mreg/_06474_ ;
wire \mreg/_06475_ ;
wire \mreg/_06476_ ;
wire \mreg/_06477_ ;
wire \mreg/_06478_ ;
wire \mreg/_06479_ ;
wire \mreg/_06480_ ;
wire \mreg/_06481_ ;
wire \mreg/_06482_ ;
wire \mreg/_06483_ ;
wire \mreg/_06484_ ;
wire \mreg/_06485_ ;
wire \mreg/_06486_ ;
wire \mreg/_06487_ ;
wire \mreg/_06488_ ;
wire \mreg/_06489_ ;
wire \mreg/_06490_ ;
wire \mreg/_06491_ ;
wire \mreg/_06492_ ;
wire \mreg/_06493_ ;
wire \mreg/_06494_ ;
wire \mreg/_06495_ ;
wire \mreg/_06496_ ;
wire \mreg/_06497_ ;
wire \mreg/_06498_ ;
wire \mreg/_06499_ ;
wire \mreg/_06500_ ;
wire \mreg/_06501_ ;
wire \mreg/_06502_ ;
wire \mreg/_06503_ ;
wire \mreg/_06504_ ;
wire \mreg/_06505_ ;
wire \mreg/_06506_ ;
wire \mreg/_06507_ ;
wire \mreg/_06508_ ;
wire \mreg/_06509_ ;
wire \mreg/_06510_ ;
wire \mreg/_06511_ ;
wire \mreg/_06512_ ;
wire \mreg/_06513_ ;
wire \mreg/_06514_ ;
wire \mreg/_06515_ ;
wire \mreg/_06516_ ;
wire \mreg/_06517_ ;
wire \mreg/_06518_ ;
wire \mreg/_06519_ ;
wire \mreg/_06520_ ;
wire \mreg/_06521_ ;
wire \mreg/_06522_ ;
wire \mreg/_06523_ ;
wire \mreg/_06524_ ;
wire \mreg/_06525_ ;
wire \mreg/_06526_ ;
wire \mreg/_06527_ ;
wire \mreg/_06528_ ;
wire \mreg/_06529_ ;
wire \mreg/_06530_ ;
wire \mreg/_06531_ ;
wire \mreg/_06532_ ;
wire \mreg/_06533_ ;
wire \mreg/_06534_ ;
wire \mreg/_06535_ ;
wire \mreg/_06536_ ;
wire \mreg/_06537_ ;
wire \mreg/_06538_ ;
wire \mreg/_06539_ ;
wire \mreg/_06540_ ;
wire \mreg/_06541_ ;
wire \mreg/_06542_ ;
wire \mreg/_06543_ ;
wire \mreg/_06544_ ;
wire \mreg/_06545_ ;
wire \mreg/_06546_ ;
wire \mreg/_06547_ ;
wire \mreg/_06548_ ;
wire \mreg/_06549_ ;
wire \mreg/_06550_ ;
wire \mreg/_06551_ ;
wire \mreg/_06552_ ;
wire \mreg/_06553_ ;
wire \mreg/_06554_ ;
wire \mreg/_06555_ ;
wire \mreg/_06556_ ;
wire \mreg/_06557_ ;
wire \mreg/_06558_ ;
wire \mreg/_06559_ ;
wire \mreg/_06560_ ;
wire \mreg/_06561_ ;
wire \mreg/_06562_ ;
wire \mreg/_06563_ ;
wire \mreg/_06564_ ;
wire \mreg/_06565_ ;
wire \mreg/_06566_ ;
wire \mreg/_06567_ ;
wire \mreg/_06568_ ;
wire \mreg/_06569_ ;
wire \mreg/_06570_ ;
wire \mreg/_06571_ ;
wire \mreg/_06572_ ;
wire \mreg/_06573_ ;
wire \mreg/_06574_ ;
wire \mreg/_06575_ ;
wire \mreg/_06576_ ;
wire \mreg/_06577_ ;
wire \mreg/_06578_ ;
wire \mreg/_06579_ ;
wire \mreg/_06580_ ;
wire \mreg/_06581_ ;
wire \mreg/_06582_ ;
wire \mreg/_06583_ ;
wire \mreg/_06584_ ;
wire \mreg/_06585_ ;
wire \mreg/_06586_ ;
wire \mreg/_06587_ ;
wire \mreg/_06588_ ;
wire \mreg/_06589_ ;
wire \mreg/_06590_ ;
wire \mreg/_06591_ ;
wire \mreg/_06592_ ;
wire \mreg/_06593_ ;
wire \mreg/_06594_ ;
wire \mreg/_06595_ ;
wire \mreg/_06596_ ;
wire \mreg/_06597_ ;
wire \mreg/_06598_ ;
wire \mreg/_06599_ ;
wire \mreg/_06600_ ;
wire \mreg/_06601_ ;
wire \mreg/_06602_ ;
wire \mreg/_06603_ ;
wire \mreg/_06604_ ;
wire \mreg/_06605_ ;
wire \mreg/_06606_ ;
wire \mreg/_06607_ ;
wire \mreg/_06608_ ;
wire \mreg/_06609_ ;
wire \mreg/_06610_ ;
wire \mreg/_06611_ ;
wire \mreg/_06612_ ;
wire \mreg/_06613_ ;
wire \mreg/_06614_ ;
wire \mreg/_06615_ ;
wire \mreg/_06616_ ;
wire \mreg/_06617_ ;
wire \mreg/_06618_ ;
wire \mreg/_06619_ ;
wire \mreg/_06620_ ;
wire \mreg/_06621_ ;
wire \mreg/_06622_ ;
wire \mreg/_06623_ ;
wire \mreg/_06624_ ;
wire \mreg/_06625_ ;
wire \mreg/_06626_ ;
wire \mreg/_06627_ ;
wire \mreg/_06628_ ;
wire \mreg/_06629_ ;
wire \mreg/_06630_ ;
wire \mreg/_06631_ ;
wire \mreg/_06632_ ;
wire \mreg/_06633_ ;
wire \mreg/_06634_ ;
wire \mreg/_06635_ ;
wire \mreg/_06636_ ;
wire \mreg/_06637_ ;
wire \mreg/_06638_ ;
wire \mreg/_06639_ ;
wire \mreg/_06640_ ;
wire \mreg/_06641_ ;
wire \mreg/_06642_ ;
wire \mreg/_06643_ ;
wire \mreg/_06644_ ;
wire \mreg/_06645_ ;
wire \mreg/_06646_ ;
wire \mreg/_06647_ ;
wire \mreg/_06648_ ;
wire \mreg/_06649_ ;
wire \mreg/_06650_ ;
wire \mreg/_06651_ ;
wire \mreg/_06652_ ;
wire \mreg/_06653_ ;
wire \mreg/_06654_ ;
wire \mreg/_06655_ ;
wire \mreg/_06656_ ;
wire \mreg/_06657_ ;
wire \mreg/_06658_ ;
wire \mreg/_06659_ ;
wire \mreg/_06660_ ;
wire \mreg/_06661_ ;
wire \mreg/_06662_ ;
wire \mreg/_06663_ ;
wire \mreg/_06664_ ;
wire \mreg/_06665_ ;
wire \mreg/_06666_ ;
wire \mreg/_06667_ ;
wire \mreg/_06668_ ;
wire \mreg/_06669_ ;
wire \mreg/_06670_ ;
wire \mreg/_06671_ ;
wire \mreg/_06672_ ;
wire \mreg/_06673_ ;
wire \mreg/_06674_ ;
wire \mreg/_06675_ ;
wire \mreg/_06676_ ;
wire \mreg/_06677_ ;
wire \mreg/_06678_ ;
wire \mreg/_06679_ ;
wire \mreg/_06680_ ;
wire \mreg/_06681_ ;
wire \mreg/_06682_ ;
wire \mreg/_06683_ ;
wire \mreg/_06684_ ;
wire \mreg/_06685_ ;
wire \mreg/_06686_ ;
wire \mreg/_06687_ ;
wire \mreg/_06688_ ;
wire \mreg/_06689_ ;
wire \mreg/_06690_ ;
wire \mreg/_06691_ ;
wire \mreg/_06692_ ;
wire \mreg/_06693_ ;
wire \mreg/_06694_ ;
wire \mreg/_06695_ ;
wire \mreg/_06696_ ;
wire \mreg/_06697_ ;
wire \mreg/_06698_ ;
wire \mreg/_06699_ ;
wire \mreg/_06700_ ;
wire \mreg/_06701_ ;
wire \mreg/_06702_ ;
wire \mreg/_06703_ ;
wire \mreg/_06704_ ;
wire \mreg/_06705_ ;
wire \mreg/_06706_ ;
wire \mreg/_06707_ ;
wire \mreg/_06708_ ;
wire \mreg/_06709_ ;
wire \mreg/_06710_ ;
wire \mreg/_06711_ ;
wire \mreg/_06712_ ;
wire \mreg/_06713_ ;
wire \mreg/_06714_ ;
wire \mreg/_06715_ ;
wire \mreg/_06716_ ;
wire \mreg/_06717_ ;
wire \mreg/_06718_ ;
wire \mreg/_06719_ ;
wire \mreg/_06720_ ;
wire \mreg/_06721_ ;
wire \mreg/_06722_ ;
wire \mreg/_06723_ ;
wire \mreg/_06724_ ;
wire \mreg/_06725_ ;
wire \mreg/_06726_ ;
wire \mreg/_06727_ ;
wire \mreg/_06728_ ;
wire \mreg/_06729_ ;
wire \mreg/_06730_ ;
wire \mreg/_06731_ ;
wire \mreg/_06732_ ;
wire \mreg/_06733_ ;
wire \mreg/_06734_ ;
wire \mreg/_06735_ ;
wire \mreg/_06736_ ;
wire \mreg/_06737_ ;
wire \mreg/_06738_ ;
wire \mreg/_06739_ ;
wire \mreg/_06740_ ;
wire \mreg/_06741_ ;
wire \mreg/_06742_ ;
wire \mreg/_06743_ ;
wire \mreg/_06744_ ;
wire \mreg/_06745_ ;
wire \mreg/_06746_ ;
wire \mreg/_06747_ ;
wire \mreg/_06748_ ;
wire \mreg/_06749_ ;
wire \mreg/_06750_ ;
wire \mreg/_06751_ ;
wire \mreg/_06752_ ;
wire \mreg/_06753_ ;
wire \mreg/_06754_ ;
wire \mreg/_06755_ ;
wire \mreg/_06756_ ;
wire \mreg/_06757_ ;
wire \mreg/_06758_ ;
wire \mreg/_06759_ ;
wire \mreg/_06760_ ;
wire \mreg/_06761_ ;
wire \mreg/_06762_ ;
wire \mreg/_06763_ ;
wire \mreg/_06764_ ;
wire \mreg/_06765_ ;
wire \mreg/_06766_ ;
wire \mreg/_06767_ ;
wire \mreg/_06768_ ;
wire \mreg/_06769_ ;
wire \mreg/_06770_ ;
wire \mreg/_06771_ ;
wire \mreg/_06772_ ;
wire \mreg/_06773_ ;
wire \mreg/_06774_ ;
wire \mreg/_06775_ ;
wire \mreg/_06776_ ;
wire \mreg/_06777_ ;
wire \mreg/_06778_ ;
wire \mreg/_06779_ ;
wire \mreg/_06780_ ;
wire \mreg/_06781_ ;
wire \mreg/_06782_ ;
wire \mreg/_06783_ ;
wire \mreg/_06784_ ;
wire \mreg/_06785_ ;
wire \mreg/_06786_ ;
wire \mreg/_06787_ ;
wire \mreg/_06788_ ;
wire \mreg/_06789_ ;
wire \mreg/_06790_ ;
wire \mreg/_06791_ ;
wire \mreg/_06792_ ;
wire \mreg/_06793_ ;
wire \mreg/_06794_ ;
wire \mreg/_06795_ ;
wire \mreg/_06796_ ;
wire \mreg/_06797_ ;
wire \mreg/_06798_ ;
wire \mreg/_06799_ ;
wire \mreg/_06800_ ;
wire \mreg/_06801_ ;
wire \mreg/_06802_ ;
wire \mreg/_06803_ ;
wire \mreg/_06804_ ;
wire \mreg/_06805_ ;
wire \mreg/_06806_ ;
wire \mreg/_06807_ ;
wire \mreg/_06808_ ;
wire \mreg/_06809_ ;
wire \mreg/_06810_ ;
wire \mreg/_06811_ ;
wire \mreg/_06812_ ;
wire \mreg/_06813_ ;
wire \mreg/_06814_ ;
wire \mreg/_06815_ ;
wire \mreg/_06816_ ;
wire \mreg/_06817_ ;
wire \mreg/_06818_ ;
wire \mreg/_06819_ ;
wire \mreg/_06820_ ;
wire \mreg/_06821_ ;
wire \mreg/_06822_ ;
wire \mreg/_06823_ ;
wire \mreg/_06824_ ;
wire \mreg/_06825_ ;
wire \mreg/_06826_ ;
wire \mreg/_06827_ ;
wire \mreg/_06828_ ;
wire \mreg/_06829_ ;
wire \mreg/_06830_ ;
wire \mreg/_06831_ ;
wire \mreg/_06832_ ;
wire \mreg/_06833_ ;
wire \mreg/_06834_ ;
wire \mreg/_06835_ ;
wire \mreg/_06836_ ;
wire \mreg/_06837_ ;
wire \mreg/_06838_ ;
wire \mreg/_06839_ ;
wire \mreg/_06840_ ;
wire \mreg/_06841_ ;
wire \mreg/_06842_ ;
wire \mreg/_06843_ ;
wire \mreg/_06844_ ;
wire \mreg/_06845_ ;
wire \mreg/_06846_ ;
wire \mreg/_06847_ ;
wire \mreg/_06848_ ;
wire \mreg/_06849_ ;
wire \mreg/_06850_ ;
wire \mreg/_06851_ ;
wire \mreg/_06852_ ;
wire \mreg/_06853_ ;
wire \mreg/_06854_ ;
wire \mreg/_06855_ ;
wire \mreg/_06856_ ;
wire \mreg/_06857_ ;
wire \mreg/_06858_ ;
wire \mreg/_06859_ ;
wire \mreg/_06860_ ;
wire \mreg/_06861_ ;
wire \mreg/_06862_ ;
wire \mreg/_06863_ ;
wire \mreg/_06864_ ;
wire \mreg/_06865_ ;
wire \mreg/_06866_ ;
wire \mreg/_06867_ ;
wire \mreg/_06868_ ;
wire \mreg/_06869_ ;
wire \mreg/_06870_ ;
wire \mreg/_06871_ ;
wire \mreg/_06872_ ;
wire \mreg/_06873_ ;
wire \mreg/_06874_ ;
wire \mreg/_06875_ ;
wire \mreg/_06876_ ;
wire \mreg/_06877_ ;
wire \mreg/_06878_ ;
wire \mreg/_06879_ ;
wire \mreg/_06880_ ;
wire \mreg/_06881_ ;
wire \mreg/_06882_ ;
wire \mreg/_06883_ ;
wire \mreg/_06884_ ;
wire \mreg/_06885_ ;
wire \mreg/_06886_ ;
wire \mreg/_06887_ ;
wire \mreg/_06888_ ;
wire \mreg/_06889_ ;
wire \mreg/_06890_ ;
wire \mreg/_06891_ ;
wire \mreg/_06892_ ;
wire \mreg/_06893_ ;
wire \mreg/_06894_ ;
wire \mreg/_06895_ ;
wire \mreg/_06896_ ;
wire \mreg/_06897_ ;
wire \mreg/_06898_ ;
wire \mreg/_06899_ ;
wire \mreg/_06900_ ;
wire \mreg/_06901_ ;
wire \mreg/_06902_ ;
wire \mreg/_06903_ ;
wire \mreg/_06904_ ;
wire \mreg/_06905_ ;
wire \mreg/_06906_ ;
wire \mreg/_06907_ ;
wire \mreg/_06908_ ;
wire \mreg/_06909_ ;
wire \mreg/_06910_ ;
wire \mreg/_06911_ ;
wire \mreg/_06912_ ;
wire \mreg/_06913_ ;
wire \mreg/_06914_ ;
wire \mreg/_06915_ ;
wire \mreg/_06916_ ;
wire \mreg/_06917_ ;
wire \mreg/_06918_ ;
wire \mreg/_06919_ ;
wire \mreg/_06920_ ;
wire \mreg/_06921_ ;
wire \mreg/_06922_ ;
wire \mreg/_06923_ ;
wire \mreg/_06924_ ;
wire \mreg/rf[10][0] ;
wire \mreg/rf[10][10] ;
wire \mreg/rf[10][11] ;
wire \mreg/rf[10][12] ;
wire \mreg/rf[10][13] ;
wire \mreg/rf[10][14] ;
wire \mreg/rf[10][15] ;
wire \mreg/rf[10][16] ;
wire \mreg/rf[10][17] ;
wire \mreg/rf[10][18] ;
wire \mreg/rf[10][19] ;
wire \mreg/rf[10][1] ;
wire \mreg/rf[10][20] ;
wire \mreg/rf[10][21] ;
wire \mreg/rf[10][22] ;
wire \mreg/rf[10][23] ;
wire \mreg/rf[10][24] ;
wire \mreg/rf[10][25] ;
wire \mreg/rf[10][26] ;
wire \mreg/rf[10][27] ;
wire \mreg/rf[10][28] ;
wire \mreg/rf[10][29] ;
wire \mreg/rf[10][2] ;
wire \mreg/rf[10][30] ;
wire \mreg/rf[10][31] ;
wire \mreg/rf[10][3] ;
wire \mreg/rf[10][4] ;
wire \mreg/rf[10][5] ;
wire \mreg/rf[10][6] ;
wire \mreg/rf[10][7] ;
wire \mreg/rf[10][8] ;
wire \mreg/rf[10][9] ;
wire \mreg/rf[11][0] ;
wire \mreg/rf[11][10] ;
wire \mreg/rf[11][11] ;
wire \mreg/rf[11][12] ;
wire \mreg/rf[11][13] ;
wire \mreg/rf[11][14] ;
wire \mreg/rf[11][15] ;
wire \mreg/rf[11][16] ;
wire \mreg/rf[11][17] ;
wire \mreg/rf[11][18] ;
wire \mreg/rf[11][19] ;
wire \mreg/rf[11][1] ;
wire \mreg/rf[11][20] ;
wire \mreg/rf[11][21] ;
wire \mreg/rf[11][22] ;
wire \mreg/rf[11][23] ;
wire \mreg/rf[11][24] ;
wire \mreg/rf[11][25] ;
wire \mreg/rf[11][26] ;
wire \mreg/rf[11][27] ;
wire \mreg/rf[11][28] ;
wire \mreg/rf[11][29] ;
wire \mreg/rf[11][2] ;
wire \mreg/rf[11][30] ;
wire \mreg/rf[11][31] ;
wire \mreg/rf[11][3] ;
wire \mreg/rf[11][4] ;
wire \mreg/rf[11][5] ;
wire \mreg/rf[11][6] ;
wire \mreg/rf[11][7] ;
wire \mreg/rf[11][8] ;
wire \mreg/rf[11][9] ;
wire \mreg/rf[12][0] ;
wire \mreg/rf[12][10] ;
wire \mreg/rf[12][11] ;
wire \mreg/rf[12][12] ;
wire \mreg/rf[12][13] ;
wire \mreg/rf[12][14] ;
wire \mreg/rf[12][15] ;
wire \mreg/rf[12][16] ;
wire \mreg/rf[12][17] ;
wire \mreg/rf[12][18] ;
wire \mreg/rf[12][19] ;
wire \mreg/rf[12][1] ;
wire \mreg/rf[12][20] ;
wire \mreg/rf[12][21] ;
wire \mreg/rf[12][22] ;
wire \mreg/rf[12][23] ;
wire \mreg/rf[12][24] ;
wire \mreg/rf[12][25] ;
wire \mreg/rf[12][26] ;
wire \mreg/rf[12][27] ;
wire \mreg/rf[12][28] ;
wire \mreg/rf[12][29] ;
wire \mreg/rf[12][2] ;
wire \mreg/rf[12][30] ;
wire \mreg/rf[12][31] ;
wire \mreg/rf[12][3] ;
wire \mreg/rf[12][4] ;
wire \mreg/rf[12][5] ;
wire \mreg/rf[12][6] ;
wire \mreg/rf[12][7] ;
wire \mreg/rf[12][8] ;
wire \mreg/rf[12][9] ;
wire \mreg/rf[13][0] ;
wire \mreg/rf[13][10] ;
wire \mreg/rf[13][11] ;
wire \mreg/rf[13][12] ;
wire \mreg/rf[13][13] ;
wire \mreg/rf[13][14] ;
wire \mreg/rf[13][15] ;
wire \mreg/rf[13][16] ;
wire \mreg/rf[13][17] ;
wire \mreg/rf[13][18] ;
wire \mreg/rf[13][19] ;
wire \mreg/rf[13][1] ;
wire \mreg/rf[13][20] ;
wire \mreg/rf[13][21] ;
wire \mreg/rf[13][22] ;
wire \mreg/rf[13][23] ;
wire \mreg/rf[13][24] ;
wire \mreg/rf[13][25] ;
wire \mreg/rf[13][26] ;
wire \mreg/rf[13][27] ;
wire \mreg/rf[13][28] ;
wire \mreg/rf[13][29] ;
wire \mreg/rf[13][2] ;
wire \mreg/rf[13][30] ;
wire \mreg/rf[13][31] ;
wire \mreg/rf[13][3] ;
wire \mreg/rf[13][4] ;
wire \mreg/rf[13][5] ;
wire \mreg/rf[13][6] ;
wire \mreg/rf[13][7] ;
wire \mreg/rf[13][8] ;
wire \mreg/rf[13][9] ;
wire \mreg/rf[14][0] ;
wire \mreg/rf[14][10] ;
wire \mreg/rf[14][11] ;
wire \mreg/rf[14][12] ;
wire \mreg/rf[14][13] ;
wire \mreg/rf[14][14] ;
wire \mreg/rf[14][15] ;
wire \mreg/rf[14][16] ;
wire \mreg/rf[14][17] ;
wire \mreg/rf[14][18] ;
wire \mreg/rf[14][19] ;
wire \mreg/rf[14][1] ;
wire \mreg/rf[14][20] ;
wire \mreg/rf[14][21] ;
wire \mreg/rf[14][22] ;
wire \mreg/rf[14][23] ;
wire \mreg/rf[14][24] ;
wire \mreg/rf[14][25] ;
wire \mreg/rf[14][26] ;
wire \mreg/rf[14][27] ;
wire \mreg/rf[14][28] ;
wire \mreg/rf[14][29] ;
wire \mreg/rf[14][2] ;
wire \mreg/rf[14][30] ;
wire \mreg/rf[14][31] ;
wire \mreg/rf[14][3] ;
wire \mreg/rf[14][4] ;
wire \mreg/rf[14][5] ;
wire \mreg/rf[14][6] ;
wire \mreg/rf[14][7] ;
wire \mreg/rf[14][8] ;
wire \mreg/rf[14][9] ;
wire \mreg/rf[15][0] ;
wire \mreg/rf[15][10] ;
wire \mreg/rf[15][11] ;
wire \mreg/rf[15][12] ;
wire \mreg/rf[15][13] ;
wire \mreg/rf[15][14] ;
wire \mreg/rf[15][15] ;
wire \mreg/rf[15][16] ;
wire \mreg/rf[15][17] ;
wire \mreg/rf[15][18] ;
wire \mreg/rf[15][19] ;
wire \mreg/rf[15][1] ;
wire \mreg/rf[15][20] ;
wire \mreg/rf[15][21] ;
wire \mreg/rf[15][22] ;
wire \mreg/rf[15][23] ;
wire \mreg/rf[15][24] ;
wire \mreg/rf[15][25] ;
wire \mreg/rf[15][26] ;
wire \mreg/rf[15][27] ;
wire \mreg/rf[15][28] ;
wire \mreg/rf[15][29] ;
wire \mreg/rf[15][2] ;
wire \mreg/rf[15][30] ;
wire \mreg/rf[15][31] ;
wire \mreg/rf[15][3] ;
wire \mreg/rf[15][4] ;
wire \mreg/rf[15][5] ;
wire \mreg/rf[15][6] ;
wire \mreg/rf[15][7] ;
wire \mreg/rf[15][8] ;
wire \mreg/rf[15][9] ;
wire \mreg/rf[16][0] ;
wire \mreg/rf[16][10] ;
wire \mreg/rf[16][11] ;
wire \mreg/rf[16][12] ;
wire \mreg/rf[16][13] ;
wire \mreg/rf[16][14] ;
wire \mreg/rf[16][15] ;
wire \mreg/rf[16][16] ;
wire \mreg/rf[16][17] ;
wire \mreg/rf[16][18] ;
wire \mreg/rf[16][19] ;
wire \mreg/rf[16][1] ;
wire \mreg/rf[16][20] ;
wire \mreg/rf[16][21] ;
wire \mreg/rf[16][22] ;
wire \mreg/rf[16][23] ;
wire \mreg/rf[16][24] ;
wire \mreg/rf[16][25] ;
wire \mreg/rf[16][26] ;
wire \mreg/rf[16][27] ;
wire \mreg/rf[16][28] ;
wire \mreg/rf[16][29] ;
wire \mreg/rf[16][2] ;
wire \mreg/rf[16][30] ;
wire \mreg/rf[16][31] ;
wire \mreg/rf[16][3] ;
wire \mreg/rf[16][4] ;
wire \mreg/rf[16][5] ;
wire \mreg/rf[16][6] ;
wire \mreg/rf[16][7] ;
wire \mreg/rf[16][8] ;
wire \mreg/rf[16][9] ;
wire \mreg/rf[17][0] ;
wire \mreg/rf[17][10] ;
wire \mreg/rf[17][11] ;
wire \mreg/rf[17][12] ;
wire \mreg/rf[17][13] ;
wire \mreg/rf[17][14] ;
wire \mreg/rf[17][15] ;
wire \mreg/rf[17][16] ;
wire \mreg/rf[17][17] ;
wire \mreg/rf[17][18] ;
wire \mreg/rf[17][19] ;
wire \mreg/rf[17][1] ;
wire \mreg/rf[17][20] ;
wire \mreg/rf[17][21] ;
wire \mreg/rf[17][22] ;
wire \mreg/rf[17][23] ;
wire \mreg/rf[17][24] ;
wire \mreg/rf[17][25] ;
wire \mreg/rf[17][26] ;
wire \mreg/rf[17][27] ;
wire \mreg/rf[17][28] ;
wire \mreg/rf[17][29] ;
wire \mreg/rf[17][2] ;
wire \mreg/rf[17][30] ;
wire \mreg/rf[17][31] ;
wire \mreg/rf[17][3] ;
wire \mreg/rf[17][4] ;
wire \mreg/rf[17][5] ;
wire \mreg/rf[17][6] ;
wire \mreg/rf[17][7] ;
wire \mreg/rf[17][8] ;
wire \mreg/rf[17][9] ;
wire \mreg/rf[18][0] ;
wire \mreg/rf[18][10] ;
wire \mreg/rf[18][11] ;
wire \mreg/rf[18][12] ;
wire \mreg/rf[18][13] ;
wire \mreg/rf[18][14] ;
wire \mreg/rf[18][15] ;
wire \mreg/rf[18][16] ;
wire \mreg/rf[18][17] ;
wire \mreg/rf[18][18] ;
wire \mreg/rf[18][19] ;
wire \mreg/rf[18][1] ;
wire \mreg/rf[18][20] ;
wire \mreg/rf[18][21] ;
wire \mreg/rf[18][22] ;
wire \mreg/rf[18][23] ;
wire \mreg/rf[18][24] ;
wire \mreg/rf[18][25] ;
wire \mreg/rf[18][26] ;
wire \mreg/rf[18][27] ;
wire \mreg/rf[18][28] ;
wire \mreg/rf[18][29] ;
wire \mreg/rf[18][2] ;
wire \mreg/rf[18][30] ;
wire \mreg/rf[18][31] ;
wire \mreg/rf[18][3] ;
wire \mreg/rf[18][4] ;
wire \mreg/rf[18][5] ;
wire \mreg/rf[18][6] ;
wire \mreg/rf[18][7] ;
wire \mreg/rf[18][8] ;
wire \mreg/rf[18][9] ;
wire \mreg/rf[19][0] ;
wire \mreg/rf[19][10] ;
wire \mreg/rf[19][11] ;
wire \mreg/rf[19][12] ;
wire \mreg/rf[19][13] ;
wire \mreg/rf[19][14] ;
wire \mreg/rf[19][15] ;
wire \mreg/rf[19][16] ;
wire \mreg/rf[19][17] ;
wire \mreg/rf[19][18] ;
wire \mreg/rf[19][19] ;
wire \mreg/rf[19][1] ;
wire \mreg/rf[19][20] ;
wire \mreg/rf[19][21] ;
wire \mreg/rf[19][22] ;
wire \mreg/rf[19][23] ;
wire \mreg/rf[19][24] ;
wire \mreg/rf[19][25] ;
wire \mreg/rf[19][26] ;
wire \mreg/rf[19][27] ;
wire \mreg/rf[19][28] ;
wire \mreg/rf[19][29] ;
wire \mreg/rf[19][2] ;
wire \mreg/rf[19][30] ;
wire \mreg/rf[19][31] ;
wire \mreg/rf[19][3] ;
wire \mreg/rf[19][4] ;
wire \mreg/rf[19][5] ;
wire \mreg/rf[19][6] ;
wire \mreg/rf[19][7] ;
wire \mreg/rf[19][8] ;
wire \mreg/rf[19][9] ;
wire \mreg/rf[1][0] ;
wire \mreg/rf[1][10] ;
wire \mreg/rf[1][11] ;
wire \mreg/rf[1][12] ;
wire \mreg/rf[1][13] ;
wire \mreg/rf[1][14] ;
wire \mreg/rf[1][15] ;
wire \mreg/rf[1][16] ;
wire \mreg/rf[1][17] ;
wire \mreg/rf[1][18] ;
wire \mreg/rf[1][19] ;
wire \mreg/rf[1][1] ;
wire \mreg/rf[1][20] ;
wire \mreg/rf[1][21] ;
wire \mreg/rf[1][22] ;
wire \mreg/rf[1][23] ;
wire \mreg/rf[1][24] ;
wire \mreg/rf[1][25] ;
wire \mreg/rf[1][26] ;
wire \mreg/rf[1][27] ;
wire \mreg/rf[1][28] ;
wire \mreg/rf[1][29] ;
wire \mreg/rf[1][2] ;
wire \mreg/rf[1][30] ;
wire \mreg/rf[1][31] ;
wire \mreg/rf[1][3] ;
wire \mreg/rf[1][4] ;
wire \mreg/rf[1][5] ;
wire \mreg/rf[1][6] ;
wire \mreg/rf[1][7] ;
wire \mreg/rf[1][8] ;
wire \mreg/rf[1][9] ;
wire \mreg/rf[20][0] ;
wire \mreg/rf[20][10] ;
wire \mreg/rf[20][11] ;
wire \mreg/rf[20][12] ;
wire \mreg/rf[20][13] ;
wire \mreg/rf[20][14] ;
wire \mreg/rf[20][15] ;
wire \mreg/rf[20][16] ;
wire \mreg/rf[20][17] ;
wire \mreg/rf[20][18] ;
wire \mreg/rf[20][19] ;
wire \mreg/rf[20][1] ;
wire \mreg/rf[20][20] ;
wire \mreg/rf[20][21] ;
wire \mreg/rf[20][22] ;
wire \mreg/rf[20][23] ;
wire \mreg/rf[20][24] ;
wire \mreg/rf[20][25] ;
wire \mreg/rf[20][26] ;
wire \mreg/rf[20][27] ;
wire \mreg/rf[20][28] ;
wire \mreg/rf[20][29] ;
wire \mreg/rf[20][2] ;
wire \mreg/rf[20][30] ;
wire \mreg/rf[20][31] ;
wire \mreg/rf[20][3] ;
wire \mreg/rf[20][4] ;
wire \mreg/rf[20][5] ;
wire \mreg/rf[20][6] ;
wire \mreg/rf[20][7] ;
wire \mreg/rf[20][8] ;
wire \mreg/rf[20][9] ;
wire \mreg/rf[21][0] ;
wire \mreg/rf[21][10] ;
wire \mreg/rf[21][11] ;
wire \mreg/rf[21][12] ;
wire \mreg/rf[21][13] ;
wire \mreg/rf[21][14] ;
wire \mreg/rf[21][15] ;
wire \mreg/rf[21][16] ;
wire \mreg/rf[21][17] ;
wire \mreg/rf[21][18] ;
wire \mreg/rf[21][19] ;
wire \mreg/rf[21][1] ;
wire \mreg/rf[21][20] ;
wire \mreg/rf[21][21] ;
wire \mreg/rf[21][22] ;
wire \mreg/rf[21][23] ;
wire \mreg/rf[21][24] ;
wire \mreg/rf[21][25] ;
wire \mreg/rf[21][26] ;
wire \mreg/rf[21][27] ;
wire \mreg/rf[21][28] ;
wire \mreg/rf[21][29] ;
wire \mreg/rf[21][2] ;
wire \mreg/rf[21][30] ;
wire \mreg/rf[21][31] ;
wire \mreg/rf[21][3] ;
wire \mreg/rf[21][4] ;
wire \mreg/rf[21][5] ;
wire \mreg/rf[21][6] ;
wire \mreg/rf[21][7] ;
wire \mreg/rf[21][8] ;
wire \mreg/rf[21][9] ;
wire \mreg/rf[22][0] ;
wire \mreg/rf[22][10] ;
wire \mreg/rf[22][11] ;
wire \mreg/rf[22][12] ;
wire \mreg/rf[22][13] ;
wire \mreg/rf[22][14] ;
wire \mreg/rf[22][15] ;
wire \mreg/rf[22][16] ;
wire \mreg/rf[22][17] ;
wire \mreg/rf[22][18] ;
wire \mreg/rf[22][19] ;
wire \mreg/rf[22][1] ;
wire \mreg/rf[22][20] ;
wire \mreg/rf[22][21] ;
wire \mreg/rf[22][22] ;
wire \mreg/rf[22][23] ;
wire \mreg/rf[22][24] ;
wire \mreg/rf[22][25] ;
wire \mreg/rf[22][26] ;
wire \mreg/rf[22][27] ;
wire \mreg/rf[22][28] ;
wire \mreg/rf[22][29] ;
wire \mreg/rf[22][2] ;
wire \mreg/rf[22][30] ;
wire \mreg/rf[22][31] ;
wire \mreg/rf[22][3] ;
wire \mreg/rf[22][4] ;
wire \mreg/rf[22][5] ;
wire \mreg/rf[22][6] ;
wire \mreg/rf[22][7] ;
wire \mreg/rf[22][8] ;
wire \mreg/rf[22][9] ;
wire \mreg/rf[23][0] ;
wire \mreg/rf[23][10] ;
wire \mreg/rf[23][11] ;
wire \mreg/rf[23][12] ;
wire \mreg/rf[23][13] ;
wire \mreg/rf[23][14] ;
wire \mreg/rf[23][15] ;
wire \mreg/rf[23][16] ;
wire \mreg/rf[23][17] ;
wire \mreg/rf[23][18] ;
wire \mreg/rf[23][19] ;
wire \mreg/rf[23][1] ;
wire \mreg/rf[23][20] ;
wire \mreg/rf[23][21] ;
wire \mreg/rf[23][22] ;
wire \mreg/rf[23][23] ;
wire \mreg/rf[23][24] ;
wire \mreg/rf[23][25] ;
wire \mreg/rf[23][26] ;
wire \mreg/rf[23][27] ;
wire \mreg/rf[23][28] ;
wire \mreg/rf[23][29] ;
wire \mreg/rf[23][2] ;
wire \mreg/rf[23][30] ;
wire \mreg/rf[23][31] ;
wire \mreg/rf[23][3] ;
wire \mreg/rf[23][4] ;
wire \mreg/rf[23][5] ;
wire \mreg/rf[23][6] ;
wire \mreg/rf[23][7] ;
wire \mreg/rf[23][8] ;
wire \mreg/rf[23][9] ;
wire \mreg/rf[24][0] ;
wire \mreg/rf[24][10] ;
wire \mreg/rf[24][11] ;
wire \mreg/rf[24][12] ;
wire \mreg/rf[24][13] ;
wire \mreg/rf[24][14] ;
wire \mreg/rf[24][15] ;
wire \mreg/rf[24][16] ;
wire \mreg/rf[24][17] ;
wire \mreg/rf[24][18] ;
wire \mreg/rf[24][19] ;
wire \mreg/rf[24][1] ;
wire \mreg/rf[24][20] ;
wire \mreg/rf[24][21] ;
wire \mreg/rf[24][22] ;
wire \mreg/rf[24][23] ;
wire \mreg/rf[24][24] ;
wire \mreg/rf[24][25] ;
wire \mreg/rf[24][26] ;
wire \mreg/rf[24][27] ;
wire \mreg/rf[24][28] ;
wire \mreg/rf[24][29] ;
wire \mreg/rf[24][2] ;
wire \mreg/rf[24][30] ;
wire \mreg/rf[24][31] ;
wire \mreg/rf[24][3] ;
wire \mreg/rf[24][4] ;
wire \mreg/rf[24][5] ;
wire \mreg/rf[24][6] ;
wire \mreg/rf[24][7] ;
wire \mreg/rf[24][8] ;
wire \mreg/rf[24][9] ;
wire \mreg/rf[25][0] ;
wire \mreg/rf[25][10] ;
wire \mreg/rf[25][11] ;
wire \mreg/rf[25][12] ;
wire \mreg/rf[25][13] ;
wire \mreg/rf[25][14] ;
wire \mreg/rf[25][15] ;
wire \mreg/rf[25][16] ;
wire \mreg/rf[25][17] ;
wire \mreg/rf[25][18] ;
wire \mreg/rf[25][19] ;
wire \mreg/rf[25][1] ;
wire \mreg/rf[25][20] ;
wire \mreg/rf[25][21] ;
wire \mreg/rf[25][22] ;
wire \mreg/rf[25][23] ;
wire \mreg/rf[25][24] ;
wire \mreg/rf[25][25] ;
wire \mreg/rf[25][26] ;
wire \mreg/rf[25][27] ;
wire \mreg/rf[25][28] ;
wire \mreg/rf[25][29] ;
wire \mreg/rf[25][2] ;
wire \mreg/rf[25][30] ;
wire \mreg/rf[25][31] ;
wire \mreg/rf[25][3] ;
wire \mreg/rf[25][4] ;
wire \mreg/rf[25][5] ;
wire \mreg/rf[25][6] ;
wire \mreg/rf[25][7] ;
wire \mreg/rf[25][8] ;
wire \mreg/rf[25][9] ;
wire \mreg/rf[26][0] ;
wire \mreg/rf[26][10] ;
wire \mreg/rf[26][11] ;
wire \mreg/rf[26][12] ;
wire \mreg/rf[26][13] ;
wire \mreg/rf[26][14] ;
wire \mreg/rf[26][15] ;
wire \mreg/rf[26][16] ;
wire \mreg/rf[26][17] ;
wire \mreg/rf[26][18] ;
wire \mreg/rf[26][19] ;
wire \mreg/rf[26][1] ;
wire \mreg/rf[26][20] ;
wire \mreg/rf[26][21] ;
wire \mreg/rf[26][22] ;
wire \mreg/rf[26][23] ;
wire \mreg/rf[26][24] ;
wire \mreg/rf[26][25] ;
wire \mreg/rf[26][26] ;
wire \mreg/rf[26][27] ;
wire \mreg/rf[26][28] ;
wire \mreg/rf[26][29] ;
wire \mreg/rf[26][2] ;
wire \mreg/rf[26][30] ;
wire \mreg/rf[26][31] ;
wire \mreg/rf[26][3] ;
wire \mreg/rf[26][4] ;
wire \mreg/rf[26][5] ;
wire \mreg/rf[26][6] ;
wire \mreg/rf[26][7] ;
wire \mreg/rf[26][8] ;
wire \mreg/rf[26][9] ;
wire \mreg/rf[27][0] ;
wire \mreg/rf[27][10] ;
wire \mreg/rf[27][11] ;
wire \mreg/rf[27][12] ;
wire \mreg/rf[27][13] ;
wire \mreg/rf[27][14] ;
wire \mreg/rf[27][15] ;
wire \mreg/rf[27][16] ;
wire \mreg/rf[27][17] ;
wire \mreg/rf[27][18] ;
wire \mreg/rf[27][19] ;
wire \mreg/rf[27][1] ;
wire \mreg/rf[27][20] ;
wire \mreg/rf[27][21] ;
wire \mreg/rf[27][22] ;
wire \mreg/rf[27][23] ;
wire \mreg/rf[27][24] ;
wire \mreg/rf[27][25] ;
wire \mreg/rf[27][26] ;
wire \mreg/rf[27][27] ;
wire \mreg/rf[27][28] ;
wire \mreg/rf[27][29] ;
wire \mreg/rf[27][2] ;
wire \mreg/rf[27][30] ;
wire \mreg/rf[27][31] ;
wire \mreg/rf[27][3] ;
wire \mreg/rf[27][4] ;
wire \mreg/rf[27][5] ;
wire \mreg/rf[27][6] ;
wire \mreg/rf[27][7] ;
wire \mreg/rf[27][8] ;
wire \mreg/rf[27][9] ;
wire \mreg/rf[28][0] ;
wire \mreg/rf[28][10] ;
wire \mreg/rf[28][11] ;
wire \mreg/rf[28][12] ;
wire \mreg/rf[28][13] ;
wire \mreg/rf[28][14] ;
wire \mreg/rf[28][15] ;
wire \mreg/rf[28][16] ;
wire \mreg/rf[28][17] ;
wire \mreg/rf[28][18] ;
wire \mreg/rf[28][19] ;
wire \mreg/rf[28][1] ;
wire \mreg/rf[28][20] ;
wire \mreg/rf[28][21] ;
wire \mreg/rf[28][22] ;
wire \mreg/rf[28][23] ;
wire \mreg/rf[28][24] ;
wire \mreg/rf[28][25] ;
wire \mreg/rf[28][26] ;
wire \mreg/rf[28][27] ;
wire \mreg/rf[28][28] ;
wire \mreg/rf[28][29] ;
wire \mreg/rf[28][2] ;
wire \mreg/rf[28][30] ;
wire \mreg/rf[28][31] ;
wire \mreg/rf[28][3] ;
wire \mreg/rf[28][4] ;
wire \mreg/rf[28][5] ;
wire \mreg/rf[28][6] ;
wire \mreg/rf[28][7] ;
wire \mreg/rf[28][8] ;
wire \mreg/rf[28][9] ;
wire \mreg/rf[29][0] ;
wire \mreg/rf[29][10] ;
wire \mreg/rf[29][11] ;
wire \mreg/rf[29][12] ;
wire \mreg/rf[29][13] ;
wire \mreg/rf[29][14] ;
wire \mreg/rf[29][15] ;
wire \mreg/rf[29][16] ;
wire \mreg/rf[29][17] ;
wire \mreg/rf[29][18] ;
wire \mreg/rf[29][19] ;
wire \mreg/rf[29][1] ;
wire \mreg/rf[29][20] ;
wire \mreg/rf[29][21] ;
wire \mreg/rf[29][22] ;
wire \mreg/rf[29][23] ;
wire \mreg/rf[29][24] ;
wire \mreg/rf[29][25] ;
wire \mreg/rf[29][26] ;
wire \mreg/rf[29][27] ;
wire \mreg/rf[29][28] ;
wire \mreg/rf[29][29] ;
wire \mreg/rf[29][2] ;
wire \mreg/rf[29][30] ;
wire \mreg/rf[29][31] ;
wire \mreg/rf[29][3] ;
wire \mreg/rf[29][4] ;
wire \mreg/rf[29][5] ;
wire \mreg/rf[29][6] ;
wire \mreg/rf[29][7] ;
wire \mreg/rf[29][8] ;
wire \mreg/rf[29][9] ;
wire \mreg/rf[2][0] ;
wire \mreg/rf[2][10] ;
wire \mreg/rf[2][11] ;
wire \mreg/rf[2][12] ;
wire \mreg/rf[2][13] ;
wire \mreg/rf[2][14] ;
wire \mreg/rf[2][15] ;
wire \mreg/rf[2][16] ;
wire \mreg/rf[2][17] ;
wire \mreg/rf[2][18] ;
wire \mreg/rf[2][19] ;
wire \mreg/rf[2][1] ;
wire \mreg/rf[2][20] ;
wire \mreg/rf[2][21] ;
wire \mreg/rf[2][22] ;
wire \mreg/rf[2][23] ;
wire \mreg/rf[2][24] ;
wire \mreg/rf[2][25] ;
wire \mreg/rf[2][26] ;
wire \mreg/rf[2][27] ;
wire \mreg/rf[2][28] ;
wire \mreg/rf[2][29] ;
wire \mreg/rf[2][2] ;
wire \mreg/rf[2][30] ;
wire \mreg/rf[2][31] ;
wire \mreg/rf[2][3] ;
wire \mreg/rf[2][4] ;
wire \mreg/rf[2][5] ;
wire \mreg/rf[2][6] ;
wire \mreg/rf[2][7] ;
wire \mreg/rf[2][8] ;
wire \mreg/rf[2][9] ;
wire \mreg/rf[30][0] ;
wire \mreg/rf[30][10] ;
wire \mreg/rf[30][11] ;
wire \mreg/rf[30][12] ;
wire \mreg/rf[30][13] ;
wire \mreg/rf[30][14] ;
wire \mreg/rf[30][15] ;
wire \mreg/rf[30][16] ;
wire \mreg/rf[30][17] ;
wire \mreg/rf[30][18] ;
wire \mreg/rf[30][19] ;
wire \mreg/rf[30][1] ;
wire \mreg/rf[30][20] ;
wire \mreg/rf[30][21] ;
wire \mreg/rf[30][22] ;
wire \mreg/rf[30][23] ;
wire \mreg/rf[30][24] ;
wire \mreg/rf[30][25] ;
wire \mreg/rf[30][26] ;
wire \mreg/rf[30][27] ;
wire \mreg/rf[30][28] ;
wire \mreg/rf[30][29] ;
wire \mreg/rf[30][2] ;
wire \mreg/rf[30][30] ;
wire \mreg/rf[30][31] ;
wire \mreg/rf[30][3] ;
wire \mreg/rf[30][4] ;
wire \mreg/rf[30][5] ;
wire \mreg/rf[30][6] ;
wire \mreg/rf[30][7] ;
wire \mreg/rf[30][8] ;
wire \mreg/rf[30][9] ;
wire \mreg/rf[31][0] ;
wire \mreg/rf[31][10] ;
wire \mreg/rf[31][11] ;
wire \mreg/rf[31][12] ;
wire \mreg/rf[31][13] ;
wire \mreg/rf[31][14] ;
wire \mreg/rf[31][15] ;
wire \mreg/rf[31][16] ;
wire \mreg/rf[31][17] ;
wire \mreg/rf[31][18] ;
wire \mreg/rf[31][19] ;
wire \mreg/rf[31][1] ;
wire \mreg/rf[31][20] ;
wire \mreg/rf[31][21] ;
wire \mreg/rf[31][22] ;
wire \mreg/rf[31][23] ;
wire \mreg/rf[31][24] ;
wire \mreg/rf[31][25] ;
wire \mreg/rf[31][26] ;
wire \mreg/rf[31][27] ;
wire \mreg/rf[31][28] ;
wire \mreg/rf[31][29] ;
wire \mreg/rf[31][2] ;
wire \mreg/rf[31][30] ;
wire \mreg/rf[31][31] ;
wire \mreg/rf[31][3] ;
wire \mreg/rf[31][4] ;
wire \mreg/rf[31][5] ;
wire \mreg/rf[31][6] ;
wire \mreg/rf[31][7] ;
wire \mreg/rf[31][8] ;
wire \mreg/rf[31][9] ;
wire \mreg/rf[3][0] ;
wire \mreg/rf[3][10] ;
wire \mreg/rf[3][11] ;
wire \mreg/rf[3][12] ;
wire \mreg/rf[3][13] ;
wire \mreg/rf[3][14] ;
wire \mreg/rf[3][15] ;
wire \mreg/rf[3][16] ;
wire \mreg/rf[3][17] ;
wire \mreg/rf[3][18] ;
wire \mreg/rf[3][19] ;
wire \mreg/rf[3][1] ;
wire \mreg/rf[3][20] ;
wire \mreg/rf[3][21] ;
wire \mreg/rf[3][22] ;
wire \mreg/rf[3][23] ;
wire \mreg/rf[3][24] ;
wire \mreg/rf[3][25] ;
wire \mreg/rf[3][26] ;
wire \mreg/rf[3][27] ;
wire \mreg/rf[3][28] ;
wire \mreg/rf[3][29] ;
wire \mreg/rf[3][2] ;
wire \mreg/rf[3][30] ;
wire \mreg/rf[3][31] ;
wire \mreg/rf[3][3] ;
wire \mreg/rf[3][4] ;
wire \mreg/rf[3][5] ;
wire \mreg/rf[3][6] ;
wire \mreg/rf[3][7] ;
wire \mreg/rf[3][8] ;
wire \mreg/rf[3][9] ;
wire \mreg/rf[4][0] ;
wire \mreg/rf[4][10] ;
wire \mreg/rf[4][11] ;
wire \mreg/rf[4][12] ;
wire \mreg/rf[4][13] ;
wire \mreg/rf[4][14] ;
wire \mreg/rf[4][15] ;
wire \mreg/rf[4][16] ;
wire \mreg/rf[4][17] ;
wire \mreg/rf[4][18] ;
wire \mreg/rf[4][19] ;
wire \mreg/rf[4][1] ;
wire \mreg/rf[4][20] ;
wire \mreg/rf[4][21] ;
wire \mreg/rf[4][22] ;
wire \mreg/rf[4][23] ;
wire \mreg/rf[4][24] ;
wire \mreg/rf[4][25] ;
wire \mreg/rf[4][26] ;
wire \mreg/rf[4][27] ;
wire \mreg/rf[4][28] ;
wire \mreg/rf[4][29] ;
wire \mreg/rf[4][2] ;
wire \mreg/rf[4][30] ;
wire \mreg/rf[4][31] ;
wire \mreg/rf[4][3] ;
wire \mreg/rf[4][4] ;
wire \mreg/rf[4][5] ;
wire \mreg/rf[4][6] ;
wire \mreg/rf[4][7] ;
wire \mreg/rf[4][8] ;
wire \mreg/rf[4][9] ;
wire \mreg/rf[5][0] ;
wire \mreg/rf[5][10] ;
wire \mreg/rf[5][11] ;
wire \mreg/rf[5][12] ;
wire \mreg/rf[5][13] ;
wire \mreg/rf[5][14] ;
wire \mreg/rf[5][15] ;
wire \mreg/rf[5][16] ;
wire \mreg/rf[5][17] ;
wire \mreg/rf[5][18] ;
wire \mreg/rf[5][19] ;
wire \mreg/rf[5][1] ;
wire \mreg/rf[5][20] ;
wire \mreg/rf[5][21] ;
wire \mreg/rf[5][22] ;
wire \mreg/rf[5][23] ;
wire \mreg/rf[5][24] ;
wire \mreg/rf[5][25] ;
wire \mreg/rf[5][26] ;
wire \mreg/rf[5][27] ;
wire \mreg/rf[5][28] ;
wire \mreg/rf[5][29] ;
wire \mreg/rf[5][2] ;
wire \mreg/rf[5][30] ;
wire \mreg/rf[5][31] ;
wire \mreg/rf[5][3] ;
wire \mreg/rf[5][4] ;
wire \mreg/rf[5][5] ;
wire \mreg/rf[5][6] ;
wire \mreg/rf[5][7] ;
wire \mreg/rf[5][8] ;
wire \mreg/rf[5][9] ;
wire \mreg/rf[6][0] ;
wire \mreg/rf[6][10] ;
wire \mreg/rf[6][11] ;
wire \mreg/rf[6][12] ;
wire \mreg/rf[6][13] ;
wire \mreg/rf[6][14] ;
wire \mreg/rf[6][15] ;
wire \mreg/rf[6][16] ;
wire \mreg/rf[6][17] ;
wire \mreg/rf[6][18] ;
wire \mreg/rf[6][19] ;
wire \mreg/rf[6][1] ;
wire \mreg/rf[6][20] ;
wire \mreg/rf[6][21] ;
wire \mreg/rf[6][22] ;
wire \mreg/rf[6][23] ;
wire \mreg/rf[6][24] ;
wire \mreg/rf[6][25] ;
wire \mreg/rf[6][26] ;
wire \mreg/rf[6][27] ;
wire \mreg/rf[6][28] ;
wire \mreg/rf[6][29] ;
wire \mreg/rf[6][2] ;
wire \mreg/rf[6][30] ;
wire \mreg/rf[6][31] ;
wire \mreg/rf[6][3] ;
wire \mreg/rf[6][4] ;
wire \mreg/rf[6][5] ;
wire \mreg/rf[6][6] ;
wire \mreg/rf[6][7] ;
wire \mreg/rf[6][8] ;
wire \mreg/rf[6][9] ;
wire \mreg/rf[7][0] ;
wire \mreg/rf[7][10] ;
wire \mreg/rf[7][11] ;
wire \mreg/rf[7][12] ;
wire \mreg/rf[7][13] ;
wire \mreg/rf[7][14] ;
wire \mreg/rf[7][15] ;
wire \mreg/rf[7][16] ;
wire \mreg/rf[7][17] ;
wire \mreg/rf[7][18] ;
wire \mreg/rf[7][19] ;
wire \mreg/rf[7][1] ;
wire \mreg/rf[7][20] ;
wire \mreg/rf[7][21] ;
wire \mreg/rf[7][22] ;
wire \mreg/rf[7][23] ;
wire \mreg/rf[7][24] ;
wire \mreg/rf[7][25] ;
wire \mreg/rf[7][26] ;
wire \mreg/rf[7][27] ;
wire \mreg/rf[7][28] ;
wire \mreg/rf[7][29] ;
wire \mreg/rf[7][2] ;
wire \mreg/rf[7][30] ;
wire \mreg/rf[7][31] ;
wire \mreg/rf[7][3] ;
wire \mreg/rf[7][4] ;
wire \mreg/rf[7][5] ;
wire \mreg/rf[7][6] ;
wire \mreg/rf[7][7] ;
wire \mreg/rf[7][8] ;
wire \mreg/rf[7][9] ;
wire \mreg/rf[8][0] ;
wire \mreg/rf[8][10] ;
wire \mreg/rf[8][11] ;
wire \mreg/rf[8][12] ;
wire \mreg/rf[8][13] ;
wire \mreg/rf[8][14] ;
wire \mreg/rf[8][15] ;
wire \mreg/rf[8][16] ;
wire \mreg/rf[8][17] ;
wire \mreg/rf[8][18] ;
wire \mreg/rf[8][19] ;
wire \mreg/rf[8][1] ;
wire \mreg/rf[8][20] ;
wire \mreg/rf[8][21] ;
wire \mreg/rf[8][22] ;
wire \mreg/rf[8][23] ;
wire \mreg/rf[8][24] ;
wire \mreg/rf[8][25] ;
wire \mreg/rf[8][26] ;
wire \mreg/rf[8][27] ;
wire \mreg/rf[8][28] ;
wire \mreg/rf[8][29] ;
wire \mreg/rf[8][2] ;
wire \mreg/rf[8][30] ;
wire \mreg/rf[8][31] ;
wire \mreg/rf[8][3] ;
wire \mreg/rf[8][4] ;
wire \mreg/rf[8][5] ;
wire \mreg/rf[8][6] ;
wire \mreg/rf[8][7] ;
wire \mreg/rf[8][8] ;
wire \mreg/rf[8][9] ;
wire \mreg/rf[9][0] ;
wire \mreg/rf[9][10] ;
wire \mreg/rf[9][11] ;
wire \mreg/rf[9][12] ;
wire \mreg/rf[9][13] ;
wire \mreg/rf[9][14] ;
wire \mreg/rf[9][15] ;
wire \mreg/rf[9][16] ;
wire \mreg/rf[9][17] ;
wire \mreg/rf[9][18] ;
wire \mreg/rf[9][19] ;
wire \mreg/rf[9][1] ;
wire \mreg/rf[9][20] ;
wire \mreg/rf[9][21] ;
wire \mreg/rf[9][22] ;
wire \mreg/rf[9][23] ;
wire \mreg/rf[9][24] ;
wire \mreg/rf[9][25] ;
wire \mreg/rf[9][26] ;
wire \mreg/rf[9][27] ;
wire \mreg/rf[9][28] ;
wire \mreg/rf[9][29] ;
wire \mreg/rf[9][2] ;
wire \mreg/rf[9][30] ;
wire \mreg/rf[9][31] ;
wire \mreg/rf[9][3] ;
wire \mreg/rf[9][4] ;
wire \mreg/rf[9][5] ;
wire \mreg/rf[9][6] ;
wire \mreg/rf[9][7] ;
wire \mreg/rf[9][8] ;
wire \mreg/rf[9][9] ;
wire \msram/_00_ ;
wire \msram/_01_ ;
wire \msram/_02_ ;
wire \msram/_03_ ;
wire \msram/_04_ ;
wire \msram/_05_ ;
wire \msram/_06_ ;
wire \msram/_07_ ;
wire \msram/_08_ ;
wire \msram/_09_ ;
wire \msram/_10_ ;
wire \msram/_11_ ;
wire \msram/_12_ ;
wire \msram/_13_ ;
wire \msram/_14_ ;

INV_X1 _352_ ( .A(_143_ ), .ZN(_196_ ) );
NOR4_X4 _353_ ( .A1(_196_ ), .A2(_144_ ), .A3(_146_ ), .A4(_145_ ), .ZN(_197_ ) );
NOR4_X4 _354_ ( .A1(_139_ ), .A2(_138_ ), .A3(_141_ ), .A4(_140_ ), .ZN(_198_ ) );
NOR4_X4 _355_ ( .A1(_152_ ), .A2(_151_ ), .A3(_155_ ), .A4(_154_ ), .ZN(_199_ ) );
NOR4_X4 _356_ ( .A1(_148_ ), .A2(_147_ ), .A3(_150_ ), .A4(_149_ ), .ZN(_200_ ) );
AND4_X2 _357_ ( .A1(_197_ ), .A2(_198_ ), .A3(_199_ ), .A4(_200_ ), .ZN(_201_ ) );
INV_X16 _358_ ( .A(_160_ ), .ZN(_202_ ) );
AND4_X1 _359_ ( .A1(_157_ ), .A2(_202_ ), .A3(_158_ ), .A4(_159_ ), .ZN(_203_ ) );
NOR2_X1 _360_ ( .A1(_156_ ), .A2(_153_ ), .ZN(_204_ ) );
AND4_X1 _361_ ( .A1(_142_ ), .A2(_203_ ), .A3(_131_ ), .A4(_204_ ), .ZN(_205_ ) );
NOR4_X1 _362_ ( .A1(_135_ ), .A2(_134_ ), .A3(_137_ ), .A4(_136_ ), .ZN(_206_ ) );
NOR4_X1 _363_ ( .A1(_162_ ), .A2(_161_ ), .A3(_133_ ), .A4(_132_ ), .ZN(_207_ ) );
AND4_X2 _364_ ( .A1(_201_ ), .A2(_205_ ), .A3(_206_ ), .A4(_207_ ), .ZN(_097_ ) );
INV_X32 _365_ ( .A(_316_ ), .ZN(_208_ ) );
NOR2_X1 _366_ ( .A1(_208_ ), .A2(_317_ ), .ZN(_209_ ) );
BUF_X4 _367_ ( .A(_209_ ), .Z(_210_ ) );
AOI22_X2 _368_ ( .A1(_210_ ), .A2(_164_ ), .B1(_317_ ), .B2(_033_ ), .ZN(_211_ ) );
INV_X1 _369_ ( .A(_317_ ), .ZN(_212_ ) );
BUF_X4 _370_ ( .A(_212_ ), .Z(_213_ ) );
BUF_X4 _371_ ( .A(_208_ ), .Z(_214_ ) );
NAND3_X1 _372_ ( .A1(_213_ ), .A2(_214_ ), .A3(_000_ ), .ZN(_215_ ) );
NAND2_X1 _373_ ( .A1(_211_ ), .A2(_215_ ), .ZN(_284_ ) );
AOI22_X1 _374_ ( .A1(_210_ ), .A2(_175_ ), .B1(_317_ ), .B2(_044_ ), .ZN(_216_ ) );
NAND3_X1 _375_ ( .A1(_213_ ), .A2(_214_ ), .A3(_011_ ), .ZN(_217_ ) );
NAND2_X1 _376_ ( .A1(_216_ ), .A2(_217_ ), .ZN(_295_ ) );
AOI22_X1 _377_ ( .A1(_210_ ), .A2(_186_ ), .B1(_317_ ), .B2(_055_ ), .ZN(_218_ ) );
NAND3_X1 _378_ ( .A1(_213_ ), .A2(_214_ ), .A3(_022_ ), .ZN(_219_ ) );
NAND2_X1 _379_ ( .A1(_218_ ), .A2(_219_ ), .ZN(_306_ ) );
AOI22_X1 _380_ ( .A1(_210_ ), .A2(_189_ ), .B1(_317_ ), .B2(_058_ ), .ZN(_220_ ) );
NAND3_X1 _381_ ( .A1(_213_ ), .A2(_214_ ), .A3(_025_ ), .ZN(_221_ ) );
NAND2_X1 _382_ ( .A1(_220_ ), .A2(_221_ ), .ZN(_309_ ) );
AOI22_X1 _383_ ( .A1(_210_ ), .A2(_190_ ), .B1(_317_ ), .B2(_059_ ), .ZN(_222_ ) );
NAND3_X1 _384_ ( .A1(_213_ ), .A2(_214_ ), .A3(_026_ ), .ZN(_223_ ) );
NAND2_X1 _385_ ( .A1(_222_ ), .A2(_223_ ), .ZN(_310_ ) );
AOI22_X1 _386_ ( .A1(_210_ ), .A2(_191_ ), .B1(_317_ ), .B2(_060_ ), .ZN(_224_ ) );
NAND3_X1 _387_ ( .A1(_213_ ), .A2(_214_ ), .A3(_027_ ), .ZN(_225_ ) );
NAND2_X1 _388_ ( .A1(_224_ ), .A2(_225_ ), .ZN(_311_ ) );
AOI22_X1 _389_ ( .A1(_210_ ), .A2(_192_ ), .B1(_317_ ), .B2(_061_ ), .ZN(_226_ ) );
NAND3_X1 _390_ ( .A1(_213_ ), .A2(_214_ ), .A3(_028_ ), .ZN(_227_ ) );
NAND2_X1 _391_ ( .A1(_226_ ), .A2(_227_ ), .ZN(_312_ ) );
AOI22_X1 _392_ ( .A1(_210_ ), .A2(_193_ ), .B1(_317_ ), .B2(_062_ ), .ZN(_228_ ) );
NAND3_X1 _393_ ( .A1(_213_ ), .A2(_214_ ), .A3(_029_ ), .ZN(_229_ ) );
NAND2_X1 _394_ ( .A1(_228_ ), .A2(_229_ ), .ZN(_313_ ) );
AOI22_X1 _395_ ( .A1(_210_ ), .A2(_194_ ), .B1(_317_ ), .B2(_063_ ), .ZN(_230_ ) );
NAND3_X1 _396_ ( .A1(_213_ ), .A2(_214_ ), .A3(_030_ ), .ZN(_231_ ) );
NAND2_X1 _397_ ( .A1(_230_ ), .A2(_231_ ), .ZN(_314_ ) );
AOI22_X1 _398_ ( .A1(_210_ ), .A2(_195_ ), .B1(_317_ ), .B2(_064_ ), .ZN(_232_ ) );
NAND3_X1 _399_ ( .A1(_213_ ), .A2(_214_ ), .A3(_031_ ), .ZN(_233_ ) );
NAND2_X1 _400_ ( .A1(_232_ ), .A2(_233_ ), .ZN(_315_ ) );
BUF_X4 _401_ ( .A(_209_ ), .Z(_234_ ) );
AOI22_X1 _402_ ( .A1(_234_ ), .A2(_165_ ), .B1(_317_ ), .B2(_034_ ), .ZN(_235_ ) );
BUF_X4 _403_ ( .A(_212_ ), .Z(_236_ ) );
BUF_X4 _404_ ( .A(_208_ ), .Z(_237_ ) );
NAND3_X1 _405_ ( .A1(_236_ ), .A2(_237_ ), .A3(_001_ ), .ZN(_238_ ) );
NAND2_X1 _406_ ( .A1(_235_ ), .A2(_238_ ), .ZN(_285_ ) );
AOI22_X1 _407_ ( .A1(_234_ ), .A2(_166_ ), .B1(_317_ ), .B2(_035_ ), .ZN(_239_ ) );
NAND3_X1 _408_ ( .A1(_236_ ), .A2(_237_ ), .A3(_002_ ), .ZN(_240_ ) );
NAND2_X1 _409_ ( .A1(_239_ ), .A2(_240_ ), .ZN(_286_ ) );
AOI22_X1 _410_ ( .A1(_234_ ), .A2(_167_ ), .B1(_317_ ), .B2(_036_ ), .ZN(_241_ ) );
NAND3_X1 _411_ ( .A1(_236_ ), .A2(_237_ ), .A3(_003_ ), .ZN(_242_ ) );
NAND2_X1 _412_ ( .A1(_241_ ), .A2(_242_ ), .ZN(_287_ ) );
AOI22_X1 _413_ ( .A1(_234_ ), .A2(_168_ ), .B1(_317_ ), .B2(_037_ ), .ZN(_243_ ) );
NAND3_X1 _414_ ( .A1(_236_ ), .A2(_237_ ), .A3(_004_ ), .ZN(_244_ ) );
NAND2_X1 _415_ ( .A1(_243_ ), .A2(_244_ ), .ZN(_288_ ) );
AOI22_X1 _416_ ( .A1(_234_ ), .A2(_169_ ), .B1(_317_ ), .B2(_038_ ), .ZN(_245_ ) );
NAND3_X1 _417_ ( .A1(_236_ ), .A2(_237_ ), .A3(_005_ ), .ZN(_246_ ) );
NAND2_X1 _418_ ( .A1(_245_ ), .A2(_246_ ), .ZN(_289_ ) );
AOI22_X1 _419_ ( .A1(_234_ ), .A2(_170_ ), .B1(_317_ ), .B2(_039_ ), .ZN(_247_ ) );
NAND3_X1 _420_ ( .A1(_236_ ), .A2(_237_ ), .A3(_006_ ), .ZN(_248_ ) );
NAND2_X1 _421_ ( .A1(_247_ ), .A2(_248_ ), .ZN(_290_ ) );
AOI22_X1 _422_ ( .A1(_234_ ), .A2(_171_ ), .B1(_317_ ), .B2(_040_ ), .ZN(_249_ ) );
NAND3_X1 _423_ ( .A1(_236_ ), .A2(_237_ ), .A3(_007_ ), .ZN(_250_ ) );
NAND2_X1 _424_ ( .A1(_249_ ), .A2(_250_ ), .ZN(_291_ ) );
AOI22_X1 _425_ ( .A1(_234_ ), .A2(_172_ ), .B1(_317_ ), .B2(_041_ ), .ZN(_251_ ) );
NAND3_X1 _426_ ( .A1(_236_ ), .A2(_237_ ), .A3(_008_ ), .ZN(_252_ ) );
NAND2_X1 _427_ ( .A1(_251_ ), .A2(_252_ ), .ZN(_292_ ) );
AOI22_X1 _428_ ( .A1(_234_ ), .A2(_173_ ), .B1(_317_ ), .B2(_042_ ), .ZN(_253_ ) );
NAND3_X1 _429_ ( .A1(_236_ ), .A2(_237_ ), .A3(_009_ ), .ZN(_254_ ) );
NAND2_X1 _430_ ( .A1(_253_ ), .A2(_254_ ), .ZN(_293_ ) );
AOI22_X1 _431_ ( .A1(_234_ ), .A2(_174_ ), .B1(_317_ ), .B2(_043_ ), .ZN(_255_ ) );
NAND3_X1 _432_ ( .A1(_236_ ), .A2(_237_ ), .A3(_010_ ), .ZN(_256_ ) );
NAND2_X1 _433_ ( .A1(_255_ ), .A2(_256_ ), .ZN(_294_ ) );
BUF_X4 _434_ ( .A(_209_ ), .Z(_257_ ) );
AOI22_X1 _435_ ( .A1(_257_ ), .A2(_176_ ), .B1(_317_ ), .B2(_045_ ), .ZN(_258_ ) );
BUF_X4 _436_ ( .A(_212_ ), .Z(_259_ ) );
BUF_X4 _437_ ( .A(_208_ ), .Z(_260_ ) );
NAND3_X1 _438_ ( .A1(_259_ ), .A2(_260_ ), .A3(_012_ ), .ZN(_261_ ) );
NAND2_X1 _439_ ( .A1(_258_ ), .A2(_261_ ), .ZN(_296_ ) );
AOI22_X1 _440_ ( .A1(_257_ ), .A2(_177_ ), .B1(_317_ ), .B2(_046_ ), .ZN(_262_ ) );
NAND3_X1 _441_ ( .A1(_259_ ), .A2(_260_ ), .A3(_013_ ), .ZN(_263_ ) );
NAND2_X1 _442_ ( .A1(_262_ ), .A2(_263_ ), .ZN(_297_ ) );
AOI22_X1 _443_ ( .A1(_257_ ), .A2(_178_ ), .B1(_317_ ), .B2(_047_ ), .ZN(_264_ ) );
NAND3_X1 _444_ ( .A1(_259_ ), .A2(_260_ ), .A3(_014_ ), .ZN(_265_ ) );
NAND2_X1 _445_ ( .A1(_264_ ), .A2(_265_ ), .ZN(_298_ ) );
AOI22_X2 _446_ ( .A1(_257_ ), .A2(_179_ ), .B1(_317_ ), .B2(_048_ ), .ZN(_266_ ) );
NAND3_X1 _447_ ( .A1(_259_ ), .A2(_260_ ), .A3(_015_ ), .ZN(_267_ ) );
NAND2_X1 _448_ ( .A1(_266_ ), .A2(_267_ ), .ZN(_299_ ) );
AOI22_X2 _449_ ( .A1(_257_ ), .A2(_180_ ), .B1(_317_ ), .B2(_049_ ), .ZN(_268_ ) );
NAND3_X1 _450_ ( .A1(_259_ ), .A2(_260_ ), .A3(_016_ ), .ZN(_269_ ) );
NAND2_X1 _451_ ( .A1(_268_ ), .A2(_269_ ), .ZN(_300_ ) );
AOI22_X2 _452_ ( .A1(_257_ ), .A2(_181_ ), .B1(_317_ ), .B2(_050_ ), .ZN(_270_ ) );
NAND3_X1 _453_ ( .A1(_259_ ), .A2(_260_ ), .A3(_017_ ), .ZN(_271_ ) );
NAND2_X1 _454_ ( .A1(_270_ ), .A2(_271_ ), .ZN(_301_ ) );
AOI22_X2 _455_ ( .A1(_257_ ), .A2(_182_ ), .B1(_317_ ), .B2(_051_ ), .ZN(_272_ ) );
NAND3_X1 _456_ ( .A1(_259_ ), .A2(_260_ ), .A3(_018_ ), .ZN(_273_ ) );
NAND2_X1 _457_ ( .A1(_272_ ), .A2(_273_ ), .ZN(_302_ ) );
AOI22_X2 _458_ ( .A1(_257_ ), .A2(_183_ ), .B1(_317_ ), .B2(_052_ ), .ZN(_274_ ) );
NAND3_X1 _459_ ( .A1(_259_ ), .A2(_260_ ), .A3(_019_ ), .ZN(_275_ ) );
NAND2_X1 _460_ ( .A1(_274_ ), .A2(_275_ ), .ZN(_303_ ) );
AOI22_X1 _461_ ( .A1(_257_ ), .A2(_184_ ), .B1(_317_ ), .B2(_053_ ), .ZN(_276_ ) );
NAND3_X1 _462_ ( .A1(_259_ ), .A2(_260_ ), .A3(_020_ ), .ZN(_277_ ) );
NAND2_X1 _463_ ( .A1(_276_ ), .A2(_277_ ), .ZN(_304_ ) );
AOI22_X1 _464_ ( .A1(_257_ ), .A2(_185_ ), .B1(_317_ ), .B2(_054_ ), .ZN(_278_ ) );
NAND3_X1 _465_ ( .A1(_259_ ), .A2(_260_ ), .A3(_021_ ), .ZN(_279_ ) );
NAND2_X1 _466_ ( .A1(_278_ ), .A2(_279_ ), .ZN(_305_ ) );
AOI22_X1 _467_ ( .A1(_209_ ), .A2(_187_ ), .B1(_317_ ), .B2(_056_ ), .ZN(_280_ ) );
NAND3_X1 _468_ ( .A1(_212_ ), .A2(_208_ ), .A3(_023_ ), .ZN(_281_ ) );
NAND2_X1 _469_ ( .A1(_280_ ), .A2(_281_ ), .ZN(_307_ ) );
AOI22_X1 _470_ ( .A1(_209_ ), .A2(_188_ ), .B1(_317_ ), .B2(_057_ ), .ZN(_282_ ) );
NAND3_X1 _471_ ( .A1(_212_ ), .A2(_208_ ), .A3(_024_ ), .ZN(_283_ ) );
NAND2_X1 _472_ ( .A1(_282_ ), .A2(_283_ ), .ZN(_308_ ) );
MUX2_X1 _473_ ( .A(_099_ ), .B(_065_ ), .S(_350_ ), .Z(_318_ ) );
MUX2_X1 _474_ ( .A(_110_ ), .B(_076_ ), .S(_350_ ), .Z(_329_ ) );
MUX2_X1 _475_ ( .A(_121_ ), .B(_087_ ), .S(_350_ ), .Z(_340_ ) );
MUX2_X1 _476_ ( .A(_124_ ), .B(_090_ ), .S(_350_ ), .Z(_343_ ) );
MUX2_X1 _477_ ( .A(_125_ ), .B(_091_ ), .S(_350_ ), .Z(_344_ ) );
MUX2_X1 _478_ ( .A(_126_ ), .B(_092_ ), .S(_350_ ), .Z(_345_ ) );
MUX2_X1 _479_ ( .A(_127_ ), .B(_093_ ), .S(_350_ ), .Z(_346_ ) );
MUX2_X1 _480_ ( .A(_128_ ), .B(_094_ ), .S(_350_ ), .Z(_347_ ) );
MUX2_X1 _481_ ( .A(_129_ ), .B(_095_ ), .S(_350_ ), .Z(_348_ ) );
MUX2_X1 _482_ ( .A(_130_ ), .B(_096_ ), .S(_350_ ), .Z(_349_ ) );
MUX2_X1 _483_ ( .A(_100_ ), .B(_066_ ), .S(_350_ ), .Z(_319_ ) );
MUX2_X1 _484_ ( .A(_101_ ), .B(_067_ ), .S(_350_ ), .Z(_320_ ) );
MUX2_X1 _485_ ( .A(_102_ ), .B(_068_ ), .S(_350_ ), .Z(_321_ ) );
MUX2_X1 _486_ ( .A(_103_ ), .B(_069_ ), .S(_350_ ), .Z(_322_ ) );
MUX2_X1 _487_ ( .A(_104_ ), .B(_070_ ), .S(_350_ ), .Z(_323_ ) );
MUX2_X1 _488_ ( .A(_105_ ), .B(_071_ ), .S(_350_ ), .Z(_324_ ) );
MUX2_X1 _489_ ( .A(_106_ ), .B(_072_ ), .S(_350_ ), .Z(_325_ ) );
MUX2_X1 _490_ ( .A(_107_ ), .B(_073_ ), .S(_350_ ), .Z(_326_ ) );
MUX2_X1 _491_ ( .A(_108_ ), .B(_074_ ), .S(_350_ ), .Z(_327_ ) );
MUX2_X1 _492_ ( .A(_109_ ), .B(_075_ ), .S(_350_ ), .Z(_328_ ) );
MUX2_X1 _493_ ( .A(_111_ ), .B(_077_ ), .S(_350_ ), .Z(_330_ ) );
MUX2_X1 _494_ ( .A(_112_ ), .B(_078_ ), .S(_350_ ), .Z(_331_ ) );
MUX2_X1 _495_ ( .A(_113_ ), .B(_079_ ), .S(_350_ ), .Z(_332_ ) );
MUX2_X1 _496_ ( .A(_114_ ), .B(_080_ ), .S(_350_ ), .Z(_333_ ) );
MUX2_X1 _497_ ( .A(_115_ ), .B(_081_ ), .S(_350_ ), .Z(_334_ ) );
MUX2_X1 _498_ ( .A(_116_ ), .B(_082_ ), .S(_350_ ), .Z(_335_ ) );
MUX2_X1 _499_ ( .A(_117_ ), .B(_083_ ), .S(_350_ ), .Z(_336_ ) );
MUX2_X1 _500_ ( .A(_118_ ), .B(_084_ ), .S(_350_ ), .Z(_337_ ) );
MUX2_X1 _501_ ( .A(_119_ ), .B(_085_ ), .S(_350_ ), .Z(_338_ ) );
MUX2_X1 _502_ ( .A(_120_ ), .B(_086_ ), .S(_350_ ), .Z(_339_ ) );
MUX2_X1 _503_ ( .A(_122_ ), .B(_088_ ), .S(_350_ ), .Z(_341_ ) );
MUX2_X1 _504_ ( .A(_123_ ), .B(_089_ ), .S(_350_ ), .Z(_342_ ) );
OR2_X1 _505_ ( .A1(_032_ ), .A2(_098_ ), .ZN(_163_ ) );
LOGIC0_X1 _506_ ( .Z(_351_ ) );
BUF_X1 _507_ ( .A(\inst[1] ), .Z(_142_ ) );
BUF_X1 _508_ ( .A(\inst[0] ), .Z(_131_ ) );
BUF_X1 _509_ ( .A(\inst[3] ), .Z(_156_ ) );
BUF_X1 _510_ ( .A(\inst[2] ), .Z(_153_ ) );
BUF_X1 _511_ ( .A(\inst[4] ), .Z(_157_ ) );
BUF_X1 _512_ ( .A(\inst[5] ), .Z(_158_ ) );
BUF_X1 _513_ ( .A(\inst[7] ), .Z(_160_ ) );
BUF_X1 _514_ ( .A(\inst[6] ), .Z(_159_ ) );
BUF_X1 _515_ ( .A(\inst[9] ), .Z(_162_ ) );
BUF_X1 _516_ ( .A(\inst[8] ), .Z(_161_ ) );
BUF_X1 _517_ ( .A(\inst[11] ), .Z(_133_ ) );
BUF_X1 _518_ ( .A(\inst[10] ), .Z(_132_ ) );
BUF_X1 _519_ ( .A(\inst[13] ), .Z(_135_ ) );
BUF_X1 _520_ ( .A(\inst[12] ), .Z(_134_ ) );
BUF_X1 _521_ ( .A(\inst[15] ), .Z(_137_ ) );
BUF_X1 _522_ ( .A(\inst[14] ), .Z(_136_ ) );
BUF_X1 _523_ ( .A(\inst[17] ), .Z(_139_ ) );
BUF_X1 _524_ ( .A(\inst[16] ), .Z(_138_ ) );
BUF_X1 _525_ ( .A(\inst[19] ), .Z(_141_ ) );
BUF_X1 _526_ ( .A(\inst[18] ), .Z(_140_ ) );
BUF_X1 _527_ ( .A(\inst[21] ), .Z(_144_ ) );
BUF_X1 _528_ ( .A(\inst[20] ), .Z(_143_ ) );
BUF_X1 _529_ ( .A(\inst[23] ), .Z(_146_ ) );
BUF_X1 _530_ ( .A(\inst[22] ), .Z(_145_ ) );
BUF_X1 _531_ ( .A(\inst[25] ), .Z(_148_ ) );
BUF_X1 _532_ ( .A(\inst[24] ), .Z(_147_ ) );
BUF_X1 _533_ ( .A(\inst[27] ), .Z(_150_ ) );
BUF_X1 _534_ ( .A(\inst[26] ), .Z(_149_ ) );
BUF_X1 _535_ ( .A(\inst[29] ), .Z(_152_ ) );
BUF_X1 _536_ ( .A(\inst[28] ), .Z(_151_ ) );
BUF_X1 _537_ ( .A(\inst[31] ), .Z(_155_ ) );
BUF_X1 _538_ ( .A(\inst[30] ), .Z(_154_ ) );
BUF_X1 _539_ ( .A(_097_ ), .Z(exit ) );
BUF_X1 _540_ ( .A(\result_ctl[1] ), .Z(_317_ ) );
BUF_X1 _541_ ( .A(\result_ctl[0] ), .Z(_316_ ) );
BUF_X1 _542_ ( .A(\csr_rdata[0] ), .Z(_033_ ) );
BUF_X1 _543_ ( .A(\mem_rdata[0] ), .Z(_164_ ) );
BUF_X1 _544_ ( .A(\alu_result[0] ), .Z(_000_ ) );
BUF_X1 _545_ ( .A(_284_ ), .Z(\result[0] ) );
BUF_X1 _546_ ( .A(\csr_rdata[1] ), .Z(_044_ ) );
BUF_X1 _547_ ( .A(\mem_rdata[1] ), .Z(_175_ ) );
BUF_X1 _548_ ( .A(\alu_result[1] ), .Z(_011_ ) );
BUF_X1 _549_ ( .A(_295_ ), .Z(\result[1] ) );
BUF_X1 _550_ ( .A(\csr_rdata[2] ), .Z(_055_ ) );
BUF_X1 _551_ ( .A(\mem_rdata[2] ), .Z(_186_ ) );
BUF_X1 _552_ ( .A(\alu_result[2] ), .Z(_022_ ) );
BUF_X1 _553_ ( .A(_306_ ), .Z(\result[2] ) );
BUF_X1 _554_ ( .A(\csr_rdata[3] ), .Z(_058_ ) );
BUF_X1 _555_ ( .A(\mem_rdata[3] ), .Z(_189_ ) );
BUF_X1 _556_ ( .A(\alu_result[3] ), .Z(_025_ ) );
BUF_X1 _557_ ( .A(_309_ ), .Z(\result[3] ) );
BUF_X1 _558_ ( .A(\csr_rdata[4] ), .Z(_059_ ) );
BUF_X1 _559_ ( .A(\mem_rdata[4] ), .Z(_190_ ) );
BUF_X1 _560_ ( .A(\alu_result[4] ), .Z(_026_ ) );
BUF_X1 _561_ ( .A(_310_ ), .Z(\result[4] ) );
BUF_X1 _562_ ( .A(\csr_rdata[5] ), .Z(_060_ ) );
BUF_X1 _563_ ( .A(\mem_rdata[5] ), .Z(_191_ ) );
BUF_X1 _564_ ( .A(\alu_result[5] ), .Z(_027_ ) );
BUF_X1 _565_ ( .A(_311_ ), .Z(\result[5] ) );
BUF_X1 _566_ ( .A(\csr_rdata[6] ), .Z(_061_ ) );
BUF_X1 _567_ ( .A(\mem_rdata[6] ), .Z(_192_ ) );
BUF_X1 _568_ ( .A(\alu_result[6] ), .Z(_028_ ) );
BUF_X1 _569_ ( .A(_312_ ), .Z(\result[6] ) );
BUF_X1 _570_ ( .A(\csr_rdata[7] ), .Z(_062_ ) );
BUF_X1 _571_ ( .A(\mem_rdata[7] ), .Z(_193_ ) );
BUF_X1 _572_ ( .A(\alu_result[7] ), .Z(_029_ ) );
BUF_X1 _573_ ( .A(_313_ ), .Z(\result[7] ) );
BUF_X1 _574_ ( .A(\csr_rdata[8] ), .Z(_063_ ) );
BUF_X1 _575_ ( .A(\mem_rdata[8] ), .Z(_194_ ) );
BUF_X1 _576_ ( .A(\alu_result[8] ), .Z(_030_ ) );
BUF_X1 _577_ ( .A(_314_ ), .Z(\result[8] ) );
BUF_X1 _578_ ( .A(\csr_rdata[9] ), .Z(_064_ ) );
BUF_X1 _579_ ( .A(\mem_rdata[9] ), .Z(_195_ ) );
BUF_X1 _580_ ( .A(\alu_result[9] ), .Z(_031_ ) );
BUF_X1 _581_ ( .A(_315_ ), .Z(\result[9] ) );
BUF_X1 _582_ ( .A(\csr_rdata[10] ), .Z(_034_ ) );
BUF_X1 _583_ ( .A(\mem_rdata[10] ), .Z(_165_ ) );
BUF_X1 _584_ ( .A(\alu_result[10] ), .Z(_001_ ) );
BUF_X1 _585_ ( .A(_285_ ), .Z(\result[10] ) );
BUF_X1 _586_ ( .A(\csr_rdata[11] ), .Z(_035_ ) );
BUF_X1 _587_ ( .A(\mem_rdata[11] ), .Z(_166_ ) );
BUF_X1 _588_ ( .A(\alu_result[11] ), .Z(_002_ ) );
BUF_X1 _589_ ( .A(_286_ ), .Z(\result[11] ) );
BUF_X1 _590_ ( .A(\csr_rdata[12] ), .Z(_036_ ) );
BUF_X1 _591_ ( .A(\mem_rdata[12] ), .Z(_167_ ) );
BUF_X1 _592_ ( .A(\alu_result[12] ), .Z(_003_ ) );
BUF_X1 _593_ ( .A(_287_ ), .Z(\result[12] ) );
BUF_X1 _594_ ( .A(\csr_rdata[13] ), .Z(_037_ ) );
BUF_X1 _595_ ( .A(\mem_rdata[13] ), .Z(_168_ ) );
BUF_X1 _596_ ( .A(\alu_result[13] ), .Z(_004_ ) );
BUF_X1 _597_ ( .A(_288_ ), .Z(\result[13] ) );
BUF_X1 _598_ ( .A(\csr_rdata[14] ), .Z(_038_ ) );
BUF_X1 _599_ ( .A(\mem_rdata[14] ), .Z(_169_ ) );
BUF_X1 _600_ ( .A(\alu_result[14] ), .Z(_005_ ) );
BUF_X1 _601_ ( .A(_289_ ), .Z(\result[14] ) );
BUF_X1 _602_ ( .A(\csr_rdata[15] ), .Z(_039_ ) );
BUF_X1 _603_ ( .A(\mem_rdata[15] ), .Z(_170_ ) );
BUF_X1 _604_ ( .A(\alu_result[15] ), .Z(_006_ ) );
BUF_X1 _605_ ( .A(_290_ ), .Z(\result[15] ) );
BUF_X1 _606_ ( .A(\csr_rdata[16] ), .Z(_040_ ) );
BUF_X1 _607_ ( .A(\mem_rdata[16] ), .Z(_171_ ) );
BUF_X1 _608_ ( .A(\alu_result[16] ), .Z(_007_ ) );
BUF_X1 _609_ ( .A(_291_ ), .Z(\result[16] ) );
BUF_X1 _610_ ( .A(\csr_rdata[17] ), .Z(_041_ ) );
BUF_X1 _611_ ( .A(\mem_rdata[17] ), .Z(_172_ ) );
BUF_X1 _612_ ( .A(\alu_result[17] ), .Z(_008_ ) );
BUF_X1 _613_ ( .A(_292_ ), .Z(\result[17] ) );
BUF_X1 _614_ ( .A(\csr_rdata[18] ), .Z(_042_ ) );
BUF_X1 _615_ ( .A(\mem_rdata[18] ), .Z(_173_ ) );
BUF_X1 _616_ ( .A(\alu_result[18] ), .Z(_009_ ) );
BUF_X1 _617_ ( .A(_293_ ), .Z(\result[18] ) );
BUF_X1 _618_ ( .A(\csr_rdata[19] ), .Z(_043_ ) );
BUF_X1 _619_ ( .A(\mem_rdata[19] ), .Z(_174_ ) );
BUF_X1 _620_ ( .A(\alu_result[19] ), .Z(_010_ ) );
BUF_X1 _621_ ( .A(_294_ ), .Z(\result[19] ) );
BUF_X1 _622_ ( .A(\csr_rdata[20] ), .Z(_045_ ) );
BUF_X1 _623_ ( .A(\mem_rdata[20] ), .Z(_176_ ) );
BUF_X1 _624_ ( .A(\alu_result[20] ), .Z(_012_ ) );
BUF_X1 _625_ ( .A(_296_ ), .Z(\result[20] ) );
BUF_X1 _626_ ( .A(\csr_rdata[21] ), .Z(_046_ ) );
BUF_X1 _627_ ( .A(\mem_rdata[21] ), .Z(_177_ ) );
BUF_X1 _628_ ( .A(\alu_result[21] ), .Z(_013_ ) );
BUF_X1 _629_ ( .A(_297_ ), .Z(\result[21] ) );
BUF_X1 _630_ ( .A(\csr_rdata[22] ), .Z(_047_ ) );
BUF_X1 _631_ ( .A(\mem_rdata[22] ), .Z(_178_ ) );
BUF_X1 _632_ ( .A(\alu_result[22] ), .Z(_014_ ) );
BUF_X1 _633_ ( .A(_298_ ), .Z(\result[22] ) );
BUF_X1 _634_ ( .A(\csr_rdata[23] ), .Z(_048_ ) );
BUF_X1 _635_ ( .A(\mem_rdata[23] ), .Z(_179_ ) );
BUF_X1 _636_ ( .A(\alu_result[23] ), .Z(_015_ ) );
BUF_X1 _637_ ( .A(_299_ ), .Z(\result[23] ) );
BUF_X1 _638_ ( .A(\csr_rdata[24] ), .Z(_049_ ) );
BUF_X1 _639_ ( .A(\mem_rdata[24] ), .Z(_180_ ) );
BUF_X1 _640_ ( .A(\alu_result[24] ), .Z(_016_ ) );
BUF_X1 _641_ ( .A(_300_ ), .Z(\result[24] ) );
BUF_X1 _642_ ( .A(\csr_rdata[25] ), .Z(_050_ ) );
BUF_X1 _643_ ( .A(\mem_rdata[25] ), .Z(_181_ ) );
BUF_X1 _644_ ( .A(\alu_result[25] ), .Z(_017_ ) );
BUF_X1 _645_ ( .A(_301_ ), .Z(\result[25] ) );
BUF_X1 _646_ ( .A(\csr_rdata[26] ), .Z(_051_ ) );
BUF_X1 _647_ ( .A(\mem_rdata[26] ), .Z(_182_ ) );
BUF_X1 _648_ ( .A(\alu_result[26] ), .Z(_018_ ) );
BUF_X1 _649_ ( .A(_302_ ), .Z(\result[26] ) );
BUF_X1 _650_ ( .A(\csr_rdata[27] ), .Z(_052_ ) );
BUF_X1 _651_ ( .A(\mem_rdata[27] ), .Z(_183_ ) );
BUF_X1 _652_ ( .A(\alu_result[27] ), .Z(_019_ ) );
BUF_X1 _653_ ( .A(_303_ ), .Z(\result[27] ) );
BUF_X1 _654_ ( .A(\csr_rdata[28] ), .Z(_053_ ) );
BUF_X1 _655_ ( .A(\mem_rdata[28] ), .Z(_184_ ) );
BUF_X1 _656_ ( .A(\alu_result[28] ), .Z(_020_ ) );
BUF_X1 _657_ ( .A(_304_ ), .Z(\result[28] ) );
BUF_X1 _658_ ( .A(\csr_rdata[29] ), .Z(_054_ ) );
BUF_X1 _659_ ( .A(\mem_rdata[29] ), .Z(_185_ ) );
BUF_X1 _660_ ( .A(\alu_result[29] ), .Z(_021_ ) );
BUF_X1 _661_ ( .A(_305_ ), .Z(\result[29] ) );
BUF_X1 _662_ ( .A(\csr_rdata[30] ), .Z(_056_ ) );
BUF_X1 _663_ ( .A(\mem_rdata[30] ), .Z(_187_ ) );
BUF_X1 _664_ ( .A(\alu_result[30] ), .Z(_023_ ) );
BUF_X1 _665_ ( .A(_307_ ), .Z(\result[30] ) );
BUF_X1 _666_ ( .A(\csr_rdata[31] ), .Z(_057_ ) );
BUF_X1 _667_ ( .A(\mem_rdata[31] ), .Z(_188_ ) );
BUF_X1 _668_ ( .A(\alu_result[31] ), .Z(_024_ ) );
BUF_X1 _669_ ( .A(_308_ ), .Z(\result[31] ) );
BUF_X1 _670_ ( .A(\exu_upc[0] ), .Z(_099_ ) );
BUF_X1 _671_ ( .A(\csr_upc[0] ), .Z(_065_ ) );
BUF_X1 _672_ ( .A(upc_ctl ), .Z(_350_ ) );
BUF_X1 _673_ ( .A(_318_ ), .Z(\upc[0] ) );
BUF_X1 _674_ ( .A(\exu_upc[1] ), .Z(_110_ ) );
BUF_X1 _675_ ( .A(\csr_upc[1] ), .Z(_076_ ) );
BUF_X1 _676_ ( .A(_329_ ), .Z(\upc[1] ) );
BUF_X1 _677_ ( .A(\exu_upc[2] ), .Z(_121_ ) );
BUF_X1 _678_ ( .A(\csr_upc[2] ), .Z(_087_ ) );
BUF_X1 _679_ ( .A(_340_ ), .Z(\upc[2] ) );
BUF_X1 _680_ ( .A(\exu_upc[3] ), .Z(_124_ ) );
BUF_X1 _681_ ( .A(\csr_upc[3] ), .Z(_090_ ) );
BUF_X1 _682_ ( .A(_343_ ), .Z(\upc[3] ) );
BUF_X1 _683_ ( .A(\exu_upc[4] ), .Z(_125_ ) );
BUF_X1 _684_ ( .A(\csr_upc[4] ), .Z(_091_ ) );
BUF_X1 _685_ ( .A(_344_ ), .Z(\upc[4] ) );
BUF_X1 _686_ ( .A(\exu_upc[5] ), .Z(_126_ ) );
BUF_X1 _687_ ( .A(\csr_upc[5] ), .Z(_092_ ) );
BUF_X1 _688_ ( .A(_345_ ), .Z(\upc[5] ) );
BUF_X1 _689_ ( .A(\exu_upc[6] ), .Z(_127_ ) );
BUF_X1 _690_ ( .A(\csr_upc[6] ), .Z(_093_ ) );
BUF_X1 _691_ ( .A(_346_ ), .Z(\upc[6] ) );
BUF_X1 _692_ ( .A(\exu_upc[7] ), .Z(_128_ ) );
BUF_X1 _693_ ( .A(\csr_upc[7] ), .Z(_094_ ) );
BUF_X1 _694_ ( .A(_347_ ), .Z(\upc[7] ) );
BUF_X1 _695_ ( .A(\exu_upc[8] ), .Z(_129_ ) );
BUF_X1 _696_ ( .A(\csr_upc[8] ), .Z(_095_ ) );
BUF_X1 _697_ ( .A(_348_ ), .Z(\upc[8] ) );
BUF_X1 _698_ ( .A(\exu_upc[9] ), .Z(_130_ ) );
BUF_X1 _699_ ( .A(\csr_upc[9] ), .Z(_096_ ) );
BUF_X1 _700_ ( .A(_349_ ), .Z(\upc[9] ) );
BUF_X1 _701_ ( .A(\exu_upc[10] ), .Z(_100_ ) );
BUF_X1 _702_ ( .A(\csr_upc[10] ), .Z(_066_ ) );
BUF_X1 _703_ ( .A(_319_ ), .Z(\upc[10] ) );
BUF_X1 _704_ ( .A(\exu_upc[11] ), .Z(_101_ ) );
BUF_X1 _705_ ( .A(\csr_upc[11] ), .Z(_067_ ) );
BUF_X1 _706_ ( .A(_320_ ), .Z(\upc[11] ) );
BUF_X1 _707_ ( .A(\exu_upc[12] ), .Z(_102_ ) );
BUF_X1 _708_ ( .A(\csr_upc[12] ), .Z(_068_ ) );
BUF_X1 _709_ ( .A(_321_ ), .Z(\upc[12] ) );
BUF_X1 _710_ ( .A(\exu_upc[13] ), .Z(_103_ ) );
BUF_X1 _711_ ( .A(\csr_upc[13] ), .Z(_069_ ) );
BUF_X1 _712_ ( .A(_322_ ), .Z(\upc[13] ) );
BUF_X1 _713_ ( .A(\exu_upc[14] ), .Z(_104_ ) );
BUF_X1 _714_ ( .A(\csr_upc[14] ), .Z(_070_ ) );
BUF_X1 _715_ ( .A(_323_ ), .Z(\upc[14] ) );
BUF_X1 _716_ ( .A(\exu_upc[15] ), .Z(_105_ ) );
BUF_X1 _717_ ( .A(\csr_upc[15] ), .Z(_071_ ) );
BUF_X1 _718_ ( .A(_324_ ), .Z(\upc[15] ) );
BUF_X1 _719_ ( .A(\exu_upc[16] ), .Z(_106_ ) );
BUF_X1 _720_ ( .A(\csr_upc[16] ), .Z(_072_ ) );
BUF_X1 _721_ ( .A(_325_ ), .Z(\upc[16] ) );
BUF_X1 _722_ ( .A(\exu_upc[17] ), .Z(_107_ ) );
BUF_X1 _723_ ( .A(\csr_upc[17] ), .Z(_073_ ) );
BUF_X1 _724_ ( .A(_326_ ), .Z(\upc[17] ) );
BUF_X1 _725_ ( .A(\exu_upc[18] ), .Z(_108_ ) );
BUF_X1 _726_ ( .A(\csr_upc[18] ), .Z(_074_ ) );
BUF_X1 _727_ ( .A(_327_ ), .Z(\upc[18] ) );
BUF_X1 _728_ ( .A(\exu_upc[19] ), .Z(_109_ ) );
BUF_X1 _729_ ( .A(\csr_upc[19] ), .Z(_075_ ) );
BUF_X1 _730_ ( .A(_328_ ), .Z(\upc[19] ) );
BUF_X1 _731_ ( .A(\exu_upc[20] ), .Z(_111_ ) );
BUF_X1 _732_ ( .A(\csr_upc[20] ), .Z(_077_ ) );
BUF_X1 _733_ ( .A(_330_ ), .Z(\upc[20] ) );
BUF_X1 _734_ ( .A(\exu_upc[21] ), .Z(_112_ ) );
BUF_X1 _735_ ( .A(\csr_upc[21] ), .Z(_078_ ) );
BUF_X1 _736_ ( .A(_331_ ), .Z(\upc[21] ) );
BUF_X1 _737_ ( .A(\exu_upc[22] ), .Z(_113_ ) );
BUF_X1 _738_ ( .A(\csr_upc[22] ), .Z(_079_ ) );
BUF_X1 _739_ ( .A(_332_ ), .Z(\upc[22] ) );
BUF_X1 _740_ ( .A(\exu_upc[23] ), .Z(_114_ ) );
BUF_X1 _741_ ( .A(\csr_upc[23] ), .Z(_080_ ) );
BUF_X1 _742_ ( .A(_333_ ), .Z(\upc[23] ) );
BUF_X1 _743_ ( .A(\exu_upc[24] ), .Z(_115_ ) );
BUF_X1 _744_ ( .A(\csr_upc[24] ), .Z(_081_ ) );
BUF_X1 _745_ ( .A(_334_ ), .Z(\upc[24] ) );
BUF_X1 _746_ ( .A(\exu_upc[25] ), .Z(_116_ ) );
BUF_X1 _747_ ( .A(\csr_upc[25] ), .Z(_082_ ) );
BUF_X1 _748_ ( .A(_335_ ), .Z(\upc[25] ) );
BUF_X1 _749_ ( .A(\exu_upc[26] ), .Z(_117_ ) );
BUF_X1 _750_ ( .A(\csr_upc[26] ), .Z(_083_ ) );
BUF_X1 _751_ ( .A(_336_ ), .Z(\upc[26] ) );
BUF_X1 _752_ ( .A(\exu_upc[27] ), .Z(_118_ ) );
BUF_X1 _753_ ( .A(\csr_upc[27] ), .Z(_084_ ) );
BUF_X1 _754_ ( .A(_337_ ), .Z(\upc[27] ) );
BUF_X1 _755_ ( .A(\exu_upc[28] ), .Z(_119_ ) );
BUF_X1 _756_ ( .A(\csr_upc[28] ), .Z(_085_ ) );
BUF_X1 _757_ ( .A(_338_ ), .Z(\upc[28] ) );
BUF_X1 _758_ ( .A(\exu_upc[29] ), .Z(_120_ ) );
BUF_X1 _759_ ( .A(\csr_upc[29] ), .Z(_086_ ) );
BUF_X1 _760_ ( .A(_339_ ), .Z(\upc[29] ) );
BUF_X1 _761_ ( .A(\exu_upc[30] ), .Z(_122_ ) );
BUF_X1 _762_ ( .A(\csr_upc[30] ), .Z(_088_ ) );
BUF_X1 _763_ ( .A(_341_ ), .Z(\upc[30] ) );
BUF_X1 _764_ ( .A(\exu_upc[31] ), .Z(_123_ ) );
BUF_X1 _765_ ( .A(\csr_upc[31] ), .Z(_089_ ) );
BUF_X1 _766_ ( .A(_342_ ), .Z(\upc[31] ) );
BUF_X1 _767_ ( .A(branch ), .Z(_032_ ) );
BUF_X1 _768_ ( .A(exu_jump ), .Z(_098_ ) );
BUF_X1 _769_ ( .A(_163_ ), .Z(jump ) );
XOR2_X1 \malu/_308_ ( .A(\malu/_307_ ), .B(\malu/_039_ ), .Z(\malu/_208_ ) );
XOR2_X1 \malu/_309_ ( .A(\malu/_307_ ), .B(\malu/_050_ ), .Z(\malu/_219_ ) );
XOR2_X1 \malu/_310_ ( .A(\malu/_307_ ), .B(\malu/_061_ ), .Z(\malu/_230_ ) );
XOR2_X1 \malu/_311_ ( .A(\malu/_307_ ), .B(\malu/_064_ ), .Z(\malu/_233_ ) );
XOR2_X1 \malu/_312_ ( .A(\malu/_307_ ), .B(\malu/_065_ ), .Z(\malu/_234_ ) );
XOR2_X1 \malu/_313_ ( .A(\malu/_307_ ), .B(\malu/_066_ ), .Z(\malu/_235_ ) );
XOR2_X1 \malu/_314_ ( .A(\malu/_307_ ), .B(\malu/_067_ ), .Z(\malu/_236_ ) );
XOR2_X1 \malu/_315_ ( .A(\malu/_307_ ), .B(\malu/_068_ ), .Z(\malu/_237_ ) );
XOR2_X1 \malu/_316_ ( .A(\malu/_307_ ), .B(\malu/_069_ ), .Z(\malu/_238_ ) );
XOR2_X1 \malu/_317_ ( .A(\malu/_307_ ), .B(\malu/_070_ ), .Z(\malu/_239_ ) );
XOR2_X1 \malu/_318_ ( .A(\malu/_307_ ), .B(\malu/_040_ ), .Z(\malu/_209_ ) );
XOR2_X1 \malu/_319_ ( .A(\malu/_307_ ), .B(\malu/_041_ ), .Z(\malu/_210_ ) );
XOR2_X1 \malu/_320_ ( .A(\malu/_307_ ), .B(\malu/_042_ ), .Z(\malu/_211_ ) );
XOR2_X1 \malu/_321_ ( .A(\malu/_307_ ), .B(\malu/_043_ ), .Z(\malu/_212_ ) );
XOR2_X1 \malu/_322_ ( .A(\malu/_307_ ), .B(\malu/_044_ ), .Z(\malu/_213_ ) );
XOR2_X1 \malu/_323_ ( .A(\malu/_307_ ), .B(\malu/_045_ ), .Z(\malu/_214_ ) );
XOR2_X1 \malu/_324_ ( .A(\malu/_307_ ), .B(\malu/_046_ ), .Z(\malu/_215_ ) );
XOR2_X1 \malu/_325_ ( .A(\malu/_307_ ), .B(\malu/_047_ ), .Z(\malu/_216_ ) );
XOR2_X1 \malu/_326_ ( .A(\malu/_307_ ), .B(\malu/_048_ ), .Z(\malu/_217_ ) );
XOR2_X1 \malu/_327_ ( .A(\malu/_307_ ), .B(\malu/_049_ ), .Z(\malu/_218_ ) );
XOR2_X1 \malu/_328_ ( .A(\malu/_307_ ), .B(\malu/_051_ ), .Z(\malu/_220_ ) );
XOR2_X1 \malu/_329_ ( .A(\malu/_307_ ), .B(\malu/_052_ ), .Z(\malu/_221_ ) );
XOR2_X1 \malu/_330_ ( .A(\malu/_307_ ), .B(\malu/_053_ ), .Z(\malu/_222_ ) );
XOR2_X1 \malu/_331_ ( .A(\malu/_307_ ), .B(\malu/_054_ ), .Z(\malu/_223_ ) );
XOR2_X1 \malu/_332_ ( .A(\malu/_307_ ), .B(\malu/_055_ ), .Z(\malu/_224_ ) );
XOR2_X1 \malu/_333_ ( .A(\malu/_307_ ), .B(\malu/_056_ ), .Z(\malu/_225_ ) );
XOR2_X1 \malu/_334_ ( .A(\malu/_307_ ), .B(\malu/_057_ ), .Z(\malu/_226_ ) );
XOR2_X1 \malu/_335_ ( .A(\malu/_307_ ), .B(\malu/_058_ ), .Z(\malu/_227_ ) );
XOR2_X1 \malu/_336_ ( .A(\malu/_307_ ), .B(\malu/_059_ ), .Z(\malu/_228_ ) );
XOR2_X1 \malu/_337_ ( .A(\malu/_307_ ), .B(\malu/_060_ ), .Z(\malu/_229_ ) );
XOR2_X1 \malu/_338_ ( .A(\malu/_307_ ), .B(\malu/_062_ ), .Z(\malu/_231_ ) );
XOR2_X1 \malu/_339_ ( .A(\malu/_307_ ), .B(\malu/_063_ ), .Z(\malu/_232_ ) );
INV_X8 \malu/_340_ ( .A(\malu/_035_ ), .ZN(\malu/_106_ ) );
INV_X32 \malu/_341_ ( .A(\malu/_038_ ), .ZN(\malu/_107_ ) );
AND4_X1 \malu/_342_ ( .A1(\malu/_106_ ), .A2(\malu/_107_ ), .A3(\malu/_036_ ), .A4(\malu/_037_ ), .ZN(\malu/_272_ ) );
INV_X32 \malu/_343_ ( .A(\malu/_037_ ), .ZN(\malu/_108_ ) );
NOR4_X1 \malu/_344_ ( .A1(\malu/_106_ ), .A2(\malu/_108_ ), .A3(\malu/_036_ ), .A4(\malu/_038_ ), .ZN(\malu/_273_ ) );
AND4_X1 \malu/_345_ ( .A1(\malu/_106_ ), .A2(\malu/_108_ ), .A3(\malu/_107_ ), .A4(\malu/_036_ ), .ZN(\malu/_072_ ) );
NOR4_X1 \malu/_346_ ( .A1(\malu/_106_ ), .A2(\malu/_036_ ), .A3(\malu/_037_ ), .A4(\malu/_038_ ), .ZN(\malu/_073_ ) );
NOR2_X4 \malu/_347_ ( .A1(\malu/_035_ ), .A2(\malu/_036_ ), .ZN(\malu/_109_ ) );
INV_X4 \malu/_348_ ( .A(\malu/_109_ ), .ZN(\malu/_110_ ) );
AOI21_X4 \malu/_349_ ( .A(\malu/_107_ ), .B1(\malu/_110_ ), .B2(\malu/_037_ ), .ZN(\malu/_111_ ) );
INV_X4 \malu/_350_ ( .A(\malu/_111_ ), .ZN(\malu/_112_ ) );
NOR2_X2 \malu/_351_ ( .A1(\malu/_037_ ), .A2(\malu/_038_ ), .ZN(\malu/_113_ ) );
NOR2_X4 \malu/_352_ ( .A1(\malu/_108_ ), .A2(\malu/_038_ ), .ZN(\malu/_114_ ) );
NAND2_X4 \malu/_353_ ( .A1(\malu/_035_ ), .A2(\malu/_036_ ), .ZN(\malu/_115_ ) );
AOI22_X4 \malu/_354_ ( .A1(\malu/_113_ ), .A2(\malu/_110_ ), .B1(\malu/_114_ ), .B2(\malu/_115_ ), .ZN(\malu/_116_ ) );
NAND3_X1 \malu/_355_ ( .A1(\malu/_112_ ), .A2(\malu/_003_ ), .A3(\malu/_116_ ), .ZN(\malu/_117_ ) );
AND3_X2 \malu/_356_ ( .A1(\malu/_110_ ), .A2(\malu/_074_ ), .A3(\malu/_113_ ), .ZN(\malu/_118_ ) );
AND2_X1 \malu/_357_ ( .A1(\malu/_114_ ), .A2(\malu/_115_ ), .ZN(\malu/_119_ ) );
AOI21_X2 \malu/_358_ ( .A(\malu/_118_ ), .B1(\malu/_274_ ), .B2(\malu/_119_ ), .ZN(\malu/_120_ ) );
XNOR2_X2 \malu/_359_ ( .A(\malu/_001_ ), .B(\malu/_027_ ), .ZN(\malu/_121_ ) );
INV_X1 \malu/_360_ ( .A(\malu/_306_ ), .ZN(\malu/_122_ ) );
OR2_X2 \malu/_361_ ( .A1(\malu/_121_ ), .A2(\malu/_122_ ), .ZN(\malu/_123_ ) );
OR2_X4 \malu/_362_ ( .A1(\malu/_000_ ), .A2(\malu/_306_ ), .ZN(\malu/_124_ ) );
AND2_X4 \malu/_363_ ( .A1(\malu/_123_ ), .A2(\malu/_124_ ), .ZN(\malu/_125_ ) );
OAI211_X2 \malu/_364_ ( .A(\malu/_117_ ), .B(\malu/_120_ ), .C1(\malu/_125_ ), .C2(\malu/_112_ ), .ZN(\malu/_240_ ) );
AND2_X4 \malu/_365_ ( .A1(\malu/_112_ ), .A2(\malu/_116_ ), .ZN(\malu/_126_ ) );
BUF_X16 \malu/_366_ ( .A(\malu/_126_ ), .Z(\malu/_127_ ) );
BUF_X4 \malu/_367_ ( .A(\malu/_119_ ), .Z(\malu/_128_ ) );
AOI22_X2 \malu/_368_ ( .A1(\malu/_127_ ), .A2(\malu/_014_ ), .B1(\malu/_285_ ), .B2(\malu/_128_ ), .ZN(\malu/_129_ ) );
CLKBUF_X1 \malu/_369_ ( .A(\malu/_110_ ), .Z(\malu/_130_ ) );
CLKBUF_X1 \malu/_370_ ( .A(\malu/_113_ ), .Z(\malu/_131_ ) );
NAND3_X1 \malu/_371_ ( .A1(\malu/_130_ ), .A2(\malu/_085_ ), .A3(\malu/_131_ ), .ZN(\malu/_132_ ) );
NAND2_X1 \malu/_372_ ( .A1(\malu/_129_ ), .A2(\malu/_132_ ), .ZN(\malu/_251_ ) );
AOI22_X2 \malu/_373_ ( .A1(\malu/_127_ ), .A2(\malu/_025_ ), .B1(\malu/_296_ ), .B2(\malu/_128_ ), .ZN(\malu/_133_ ) );
NAND3_X1 \malu/_374_ ( .A1(\malu/_130_ ), .A2(\malu/_096_ ), .A3(\malu/_131_ ), .ZN(\malu/_134_ ) );
NAND2_X1 \malu/_375_ ( .A1(\malu/_133_ ), .A2(\malu/_134_ ), .ZN(\malu/_262_ ) );
AOI22_X2 \malu/_376_ ( .A1(\malu/_127_ ), .A2(\malu/_028_ ), .B1(\malu/_299_ ), .B2(\malu/_128_ ), .ZN(\malu/_135_ ) );
NAND3_X1 \malu/_377_ ( .A1(\malu/_130_ ), .A2(\malu/_099_ ), .A3(\malu/_131_ ), .ZN(\malu/_136_ ) );
NAND2_X1 \malu/_378_ ( .A1(\malu/_135_ ), .A2(\malu/_136_ ), .ZN(\malu/_265_ ) );
AOI22_X2 \malu/_379_ ( .A1(\malu/_127_ ), .A2(\malu/_029_ ), .B1(\malu/_300_ ), .B2(\malu/_128_ ), .ZN(\malu/_137_ ) );
NAND3_X1 \malu/_380_ ( .A1(\malu/_130_ ), .A2(\malu/_100_ ), .A3(\malu/_131_ ), .ZN(\malu/_138_ ) );
NAND2_X1 \malu/_381_ ( .A1(\malu/_137_ ), .A2(\malu/_138_ ), .ZN(\malu/_266_ ) );
AOI22_X2 \malu/_382_ ( .A1(\malu/_127_ ), .A2(\malu/_030_ ), .B1(\malu/_301_ ), .B2(\malu/_128_ ), .ZN(\malu/_139_ ) );
NAND3_X1 \malu/_383_ ( .A1(\malu/_130_ ), .A2(\malu/_101_ ), .A3(\malu/_131_ ), .ZN(\malu/_140_ ) );
NAND2_X1 \malu/_384_ ( .A1(\malu/_139_ ), .A2(\malu/_140_ ), .ZN(\malu/_267_ ) );
AOI22_X2 \malu/_385_ ( .A1(\malu/_127_ ), .A2(\malu/_031_ ), .B1(\malu/_302_ ), .B2(\malu/_128_ ), .ZN(\malu/_141_ ) );
NAND3_X1 \malu/_386_ ( .A1(\malu/_130_ ), .A2(\malu/_102_ ), .A3(\malu/_131_ ), .ZN(\malu/_142_ ) );
NAND2_X1 \malu/_387_ ( .A1(\malu/_141_ ), .A2(\malu/_142_ ), .ZN(\malu/_268_ ) );
AOI22_X2 \malu/_388_ ( .A1(\malu/_127_ ), .A2(\malu/_032_ ), .B1(\malu/_303_ ), .B2(\malu/_128_ ), .ZN(\malu/_143_ ) );
NAND3_X1 \malu/_389_ ( .A1(\malu/_130_ ), .A2(\malu/_103_ ), .A3(\malu/_131_ ), .ZN(\malu/_144_ ) );
NAND2_X1 \malu/_390_ ( .A1(\malu/_143_ ), .A2(\malu/_144_ ), .ZN(\malu/_269_ ) );
AOI22_X2 \malu/_391_ ( .A1(\malu/_127_ ), .A2(\malu/_033_ ), .B1(\malu/_304_ ), .B2(\malu/_128_ ), .ZN(\malu/_145_ ) );
NAND3_X1 \malu/_392_ ( .A1(\malu/_130_ ), .A2(\malu/_104_ ), .A3(\malu/_131_ ), .ZN(\malu/_146_ ) );
NAND2_X1 \malu/_393_ ( .A1(\malu/_145_ ), .A2(\malu/_146_ ), .ZN(\malu/_270_ ) );
AOI22_X2 \malu/_394_ ( .A1(\malu/_127_ ), .A2(\malu/_034_ ), .B1(\malu/_305_ ), .B2(\malu/_128_ ), .ZN(\malu/_147_ ) );
NAND3_X1 \malu/_395_ ( .A1(\malu/_130_ ), .A2(\malu/_105_ ), .A3(\malu/_131_ ), .ZN(\malu/_148_ ) );
NAND2_X1 \malu/_396_ ( .A1(\malu/_147_ ), .A2(\malu/_148_ ), .ZN(\malu/_271_ ) );
AOI22_X2 \malu/_397_ ( .A1(\malu/_127_ ), .A2(\malu/_004_ ), .B1(\malu/_275_ ), .B2(\malu/_128_ ), .ZN(\malu/_149_ ) );
NAND3_X1 \malu/_398_ ( .A1(\malu/_130_ ), .A2(\malu/_075_ ), .A3(\malu/_131_ ), .ZN(\malu/_150_ ) );
NAND2_X1 \malu/_399_ ( .A1(\malu/_149_ ), .A2(\malu/_150_ ), .ZN(\malu/_241_ ) );
BUF_X16 \malu/_400_ ( .A(\malu/_126_ ), .Z(\malu/_151_ ) );
BUF_X4 \malu/_401_ ( .A(\malu/_119_ ), .Z(\malu/_152_ ) );
AOI22_X2 \malu/_402_ ( .A1(\malu/_151_ ), .A2(\malu/_005_ ), .B1(\malu/_276_ ), .B2(\malu/_152_ ), .ZN(\malu/_153_ ) );
CLKBUF_X1 \malu/_403_ ( .A(\malu/_110_ ), .Z(\malu/_154_ ) );
CLKBUF_X1 \malu/_404_ ( .A(\malu/_113_ ), .Z(\malu/_155_ ) );
NAND3_X1 \malu/_405_ ( .A1(\malu/_154_ ), .A2(\malu/_076_ ), .A3(\malu/_155_ ), .ZN(\malu/_156_ ) );
NAND2_X1 \malu/_406_ ( .A1(\malu/_153_ ), .A2(\malu/_156_ ), .ZN(\malu/_242_ ) );
AOI22_X2 \malu/_407_ ( .A1(\malu/_151_ ), .A2(\malu/_006_ ), .B1(\malu/_277_ ), .B2(\malu/_152_ ), .ZN(\malu/_157_ ) );
NAND3_X1 \malu/_408_ ( .A1(\malu/_154_ ), .A2(\malu/_077_ ), .A3(\malu/_155_ ), .ZN(\malu/_158_ ) );
NAND2_X1 \malu/_409_ ( .A1(\malu/_157_ ), .A2(\malu/_158_ ), .ZN(\malu/_243_ ) );
AOI22_X2 \malu/_410_ ( .A1(\malu/_151_ ), .A2(\malu/_007_ ), .B1(\malu/_278_ ), .B2(\malu/_152_ ), .ZN(\malu/_159_ ) );
NAND3_X1 \malu/_411_ ( .A1(\malu/_154_ ), .A2(\malu/_078_ ), .A3(\malu/_155_ ), .ZN(\malu/_160_ ) );
NAND2_X1 \malu/_412_ ( .A1(\malu/_159_ ), .A2(\malu/_160_ ), .ZN(\malu/_244_ ) );
AOI22_X2 \malu/_413_ ( .A1(\malu/_151_ ), .A2(\malu/_008_ ), .B1(\malu/_279_ ), .B2(\malu/_152_ ), .ZN(\malu/_161_ ) );
NAND3_X1 \malu/_414_ ( .A1(\malu/_154_ ), .A2(\malu/_079_ ), .A3(\malu/_155_ ), .ZN(\malu/_162_ ) );
NAND2_X1 \malu/_415_ ( .A1(\malu/_161_ ), .A2(\malu/_162_ ), .ZN(\malu/_245_ ) );
AOI22_X2 \malu/_416_ ( .A1(\malu/_151_ ), .A2(\malu/_009_ ), .B1(\malu/_280_ ), .B2(\malu/_152_ ), .ZN(\malu/_163_ ) );
NAND3_X1 \malu/_417_ ( .A1(\malu/_154_ ), .A2(\malu/_080_ ), .A3(\malu/_155_ ), .ZN(\malu/_164_ ) );
NAND2_X1 \malu/_418_ ( .A1(\malu/_163_ ), .A2(\malu/_164_ ), .ZN(\malu/_246_ ) );
AOI22_X2 \malu/_419_ ( .A1(\malu/_151_ ), .A2(\malu/_010_ ), .B1(\malu/_281_ ), .B2(\malu/_152_ ), .ZN(\malu/_165_ ) );
NAND3_X1 \malu/_420_ ( .A1(\malu/_154_ ), .A2(\malu/_081_ ), .A3(\malu/_155_ ), .ZN(\malu/_166_ ) );
NAND2_X1 \malu/_421_ ( .A1(\malu/_165_ ), .A2(\malu/_166_ ), .ZN(\malu/_247_ ) );
AOI22_X2 \malu/_422_ ( .A1(\malu/_151_ ), .A2(\malu/_011_ ), .B1(\malu/_282_ ), .B2(\malu/_152_ ), .ZN(\malu/_167_ ) );
NAND3_X1 \malu/_423_ ( .A1(\malu/_154_ ), .A2(\malu/_082_ ), .A3(\malu/_155_ ), .ZN(\malu/_168_ ) );
NAND2_X1 \malu/_424_ ( .A1(\malu/_167_ ), .A2(\malu/_168_ ), .ZN(\malu/_248_ ) );
AOI22_X2 \malu/_425_ ( .A1(\malu/_151_ ), .A2(\malu/_012_ ), .B1(\malu/_283_ ), .B2(\malu/_152_ ), .ZN(\malu/_169_ ) );
NAND3_X1 \malu/_426_ ( .A1(\malu/_154_ ), .A2(\malu/_083_ ), .A3(\malu/_155_ ), .ZN(\malu/_170_ ) );
NAND2_X1 \malu/_427_ ( .A1(\malu/_169_ ), .A2(\malu/_170_ ), .ZN(\malu/_249_ ) );
AOI22_X2 \malu/_428_ ( .A1(\malu/_151_ ), .A2(\malu/_013_ ), .B1(\malu/_284_ ), .B2(\malu/_152_ ), .ZN(\malu/_171_ ) );
NAND3_X1 \malu/_429_ ( .A1(\malu/_154_ ), .A2(\malu/_084_ ), .A3(\malu/_155_ ), .ZN(\malu/_172_ ) );
NAND2_X1 \malu/_430_ ( .A1(\malu/_171_ ), .A2(\malu/_172_ ), .ZN(\malu/_250_ ) );
AOI22_X2 \malu/_431_ ( .A1(\malu/_151_ ), .A2(\malu/_015_ ), .B1(\malu/_286_ ), .B2(\malu/_152_ ), .ZN(\malu/_173_ ) );
NAND3_X1 \malu/_432_ ( .A1(\malu/_154_ ), .A2(\malu/_086_ ), .A3(\malu/_155_ ), .ZN(\malu/_174_ ) );
NAND2_X1 \malu/_433_ ( .A1(\malu/_173_ ), .A2(\malu/_174_ ), .ZN(\malu/_252_ ) );
BUF_X16 \malu/_434_ ( .A(\malu/_126_ ), .Z(\malu/_175_ ) );
BUF_X4 \malu/_435_ ( .A(\malu/_119_ ), .Z(\malu/_176_ ) );
AOI22_X2 \malu/_436_ ( .A1(\malu/_175_ ), .A2(\malu/_016_ ), .B1(\malu/_287_ ), .B2(\malu/_176_ ), .ZN(\malu/_177_ ) );
CLKBUF_X1 \malu/_437_ ( .A(\malu/_110_ ), .Z(\malu/_178_ ) );
CLKBUF_X1 \malu/_438_ ( .A(\malu/_113_ ), .Z(\malu/_179_ ) );
NAND3_X1 \malu/_439_ ( .A1(\malu/_178_ ), .A2(\malu/_087_ ), .A3(\malu/_179_ ), .ZN(\malu/_180_ ) );
NAND2_X1 \malu/_440_ ( .A1(\malu/_177_ ), .A2(\malu/_180_ ), .ZN(\malu/_253_ ) );
AOI22_X2 \malu/_441_ ( .A1(\malu/_175_ ), .A2(\malu/_017_ ), .B1(\malu/_288_ ), .B2(\malu/_176_ ), .ZN(\malu/_181_ ) );
NAND3_X1 \malu/_442_ ( .A1(\malu/_178_ ), .A2(\malu/_088_ ), .A3(\malu/_179_ ), .ZN(\malu/_182_ ) );
NAND2_X1 \malu/_443_ ( .A1(\malu/_181_ ), .A2(\malu/_182_ ), .ZN(\malu/_254_ ) );
AOI22_X2 \malu/_444_ ( .A1(\malu/_175_ ), .A2(\malu/_018_ ), .B1(\malu/_289_ ), .B2(\malu/_176_ ), .ZN(\malu/_183_ ) );
NAND3_X1 \malu/_445_ ( .A1(\malu/_178_ ), .A2(\malu/_089_ ), .A3(\malu/_179_ ), .ZN(\malu/_184_ ) );
NAND2_X1 \malu/_446_ ( .A1(\malu/_183_ ), .A2(\malu/_184_ ), .ZN(\malu/_255_ ) );
AOI22_X2 \malu/_447_ ( .A1(\malu/_175_ ), .A2(\malu/_019_ ), .B1(\malu/_290_ ), .B2(\malu/_176_ ), .ZN(\malu/_185_ ) );
NAND3_X1 \malu/_448_ ( .A1(\malu/_178_ ), .A2(\malu/_090_ ), .A3(\malu/_179_ ), .ZN(\malu/_186_ ) );
NAND2_X1 \malu/_449_ ( .A1(\malu/_185_ ), .A2(\malu/_186_ ), .ZN(\malu/_256_ ) );
AOI22_X2 \malu/_450_ ( .A1(\malu/_175_ ), .A2(\malu/_020_ ), .B1(\malu/_291_ ), .B2(\malu/_176_ ), .ZN(\malu/_187_ ) );
NAND3_X1 \malu/_451_ ( .A1(\malu/_178_ ), .A2(\malu/_091_ ), .A3(\malu/_179_ ), .ZN(\malu/_188_ ) );
NAND2_X1 \malu/_452_ ( .A1(\malu/_187_ ), .A2(\malu/_188_ ), .ZN(\malu/_257_ ) );
AOI22_X2 \malu/_453_ ( .A1(\malu/_175_ ), .A2(\malu/_021_ ), .B1(\malu/_292_ ), .B2(\malu/_176_ ), .ZN(\malu/_189_ ) );
NAND3_X1 \malu/_454_ ( .A1(\malu/_178_ ), .A2(\malu/_092_ ), .A3(\malu/_179_ ), .ZN(\malu/_190_ ) );
NAND2_X1 \malu/_455_ ( .A1(\malu/_189_ ), .A2(\malu/_190_ ), .ZN(\malu/_258_ ) );
AOI22_X2 \malu/_456_ ( .A1(\malu/_175_ ), .A2(\malu/_022_ ), .B1(\malu/_293_ ), .B2(\malu/_176_ ), .ZN(\malu/_191_ ) );
NAND3_X1 \malu/_457_ ( .A1(\malu/_178_ ), .A2(\malu/_093_ ), .A3(\malu/_179_ ), .ZN(\malu/_192_ ) );
NAND2_X1 \malu/_458_ ( .A1(\malu/_191_ ), .A2(\malu/_192_ ), .ZN(\malu/_259_ ) );
AOI22_X2 \malu/_459_ ( .A1(\malu/_175_ ), .A2(\malu/_023_ ), .B1(\malu/_294_ ), .B2(\malu/_176_ ), .ZN(\malu/_193_ ) );
NAND3_X1 \malu/_460_ ( .A1(\malu/_178_ ), .A2(\malu/_094_ ), .A3(\malu/_179_ ), .ZN(\malu/_194_ ) );
NAND2_X1 \malu/_461_ ( .A1(\malu/_193_ ), .A2(\malu/_194_ ), .ZN(\malu/_260_ ) );
AOI22_X2 \malu/_462_ ( .A1(\malu/_175_ ), .A2(\malu/_024_ ), .B1(\malu/_295_ ), .B2(\malu/_176_ ), .ZN(\malu/_195_ ) );
NAND3_X1 \malu/_463_ ( .A1(\malu/_178_ ), .A2(\malu/_095_ ), .A3(\malu/_179_ ), .ZN(\malu/_196_ ) );
NAND2_X1 \malu/_464_ ( .A1(\malu/_195_ ), .A2(\malu/_196_ ), .ZN(\malu/_261_ ) );
AOI22_X2 \malu/_465_ ( .A1(\malu/_175_ ), .A2(\malu/_026_ ), .B1(\malu/_297_ ), .B2(\malu/_176_ ), .ZN(\malu/_197_ ) );
NAND3_X1 \malu/_466_ ( .A1(\malu/_178_ ), .A2(\malu/_097_ ), .A3(\malu/_179_ ), .ZN(\malu/_198_ ) );
NAND2_X1 \malu/_467_ ( .A1(\malu/_197_ ), .A2(\malu/_198_ ), .ZN(\malu/_263_ ) );
AOI22_X1 \malu/_468_ ( .A1(\malu/_126_ ), .A2(\malu/_027_ ), .B1(\malu/_298_ ), .B2(\malu/_119_ ), .ZN(\malu/_199_ ) );
NAND3_X1 \malu/_469_ ( .A1(\malu/_110_ ), .A2(\malu/_098_ ), .A3(\malu/_113_ ), .ZN(\malu/_200_ ) );
NAND2_X1 \malu/_470_ ( .A1(\malu/_199_ ), .A2(\malu/_200_ ), .ZN(\malu/_264_ ) );
NAND2_X1 \malu/_471_ ( .A1(\malu/_106_ ), .A2(\malu/_036_ ), .ZN(\malu/_201_ ) );
NAND2_X1 \malu/_472_ ( .A1(\malu/_108_ ), .A2(\malu/_038_ ), .ZN(\malu/_202_ ) );
OR3_X2 \malu/_473_ ( .A1(\malu/_125_ ), .A2(\malu/_201_ ), .A3(\malu/_202_ ), .ZN(\malu/_203_ ) );
OR4_X1 \malu/_474_ ( .A1(\malu/_106_ ), .A2(\malu/_202_ ), .A3(\malu/_036_ ), .A4(\malu/_002_ ), .ZN(\malu/_204_ ) );
NAND4_X1 \malu/_475_ ( .A1(\malu/_109_ ), .A2(\malu/_108_ ), .A3(\malu/_038_ ), .A4(\malu/_002_ ), .ZN(\malu/_205_ ) );
NOR3_X1 \malu/_476_ ( .A1(\malu/_115_ ), .A2(\malu/_107_ ), .A3(\malu/_037_ ), .ZN(\malu/_206_ ) );
OAI211_X2 \malu/_477_ ( .A(\malu/_206_ ), .B(\malu/_124_ ), .C1(\malu/_121_ ), .C2(\malu/_122_ ), .ZN(\malu/_207_ ) );
NAND4_X1 \malu/_478_ ( .A1(\malu/_203_ ), .A2(\malu/_204_ ), .A3(\malu/_205_ ), .A4(\malu/_207_ ), .ZN(\malu/_071_ ) );
BUF_X1 \malu/_479_ ( .A(alu_sub ), .Z(\malu/_307_ ) );
BUF_X1 \malu/_480_ ( .A(\alu_b[0] ), .Z(\malu/_039_ ) );
BUF_X1 \malu/_481_ ( .A(\malu/_208_ ), .Z(\malu/r[0] ) );
BUF_X1 \malu/_482_ ( .A(\alu_b[1] ), .Z(\malu/_050_ ) );
BUF_X1 \malu/_483_ ( .A(\malu/_219_ ), .Z(\malu/r[1] ) );
BUF_X1 \malu/_484_ ( .A(\alu_b[2] ), .Z(\malu/_061_ ) );
BUF_X1 \malu/_485_ ( .A(\malu/_230_ ), .Z(\malu/r[2] ) );
BUF_X1 \malu/_486_ ( .A(\alu_b[3] ), .Z(\malu/_064_ ) );
BUF_X1 \malu/_487_ ( .A(\malu/_233_ ), .Z(\malu/r[3] ) );
BUF_X1 \malu/_488_ ( .A(\alu_b[4] ), .Z(\malu/_065_ ) );
BUF_X1 \malu/_489_ ( .A(\malu/_234_ ), .Z(\malu/r[4] ) );
BUF_X1 \malu/_490_ ( .A(\alu_b[5] ), .Z(\malu/_066_ ) );
BUF_X1 \malu/_491_ ( .A(\malu/_235_ ), .Z(\malu/r[5] ) );
BUF_X1 \malu/_492_ ( .A(\alu_b[6] ), .Z(\malu/_067_ ) );
BUF_X1 \malu/_493_ ( .A(\malu/_236_ ), .Z(\malu/r[6] ) );
BUF_X1 \malu/_494_ ( .A(\alu_b[7] ), .Z(\malu/_068_ ) );
BUF_X1 \malu/_495_ ( .A(\malu/_237_ ), .Z(\malu/r[7] ) );
BUF_X1 \malu/_496_ ( .A(\alu_b[8] ), .Z(\malu/_069_ ) );
BUF_X1 \malu/_497_ ( .A(\malu/_238_ ), .Z(\malu/r[8] ) );
BUF_X1 \malu/_498_ ( .A(\alu_b[9] ), .Z(\malu/_070_ ) );
BUF_X1 \malu/_499_ ( .A(\malu/_239_ ), .Z(\malu/r[9] ) );
BUF_X1 \malu/_500_ ( .A(\alu_b[10] ), .Z(\malu/_040_ ) );
BUF_X1 \malu/_501_ ( .A(\malu/_209_ ), .Z(\malu/r[10] ) );
BUF_X1 \malu/_502_ ( .A(\alu_b[11] ), .Z(\malu/_041_ ) );
BUF_X1 \malu/_503_ ( .A(\malu/_210_ ), .Z(\malu/r[11] ) );
BUF_X1 \malu/_504_ ( .A(\alu_b[12] ), .Z(\malu/_042_ ) );
BUF_X1 \malu/_505_ ( .A(\malu/_211_ ), .Z(\malu/r[12] ) );
BUF_X1 \malu/_506_ ( .A(\alu_b[13] ), .Z(\malu/_043_ ) );
BUF_X1 \malu/_507_ ( .A(\malu/_212_ ), .Z(\malu/r[13] ) );
BUF_X1 \malu/_508_ ( .A(\alu_b[14] ), .Z(\malu/_044_ ) );
BUF_X1 \malu/_509_ ( .A(\malu/_213_ ), .Z(\malu/r[14] ) );
BUF_X1 \malu/_510_ ( .A(\alu_b[15] ), .Z(\malu/_045_ ) );
BUF_X1 \malu/_511_ ( .A(\malu/_214_ ), .Z(\malu/r[15] ) );
BUF_X1 \malu/_512_ ( .A(\alu_b[16] ), .Z(\malu/_046_ ) );
BUF_X1 \malu/_513_ ( .A(\malu/_215_ ), .Z(\malu/r[16] ) );
BUF_X1 \malu/_514_ ( .A(\alu_b[17] ), .Z(\malu/_047_ ) );
BUF_X1 \malu/_515_ ( .A(\malu/_216_ ), .Z(\malu/r[17] ) );
BUF_X1 \malu/_516_ ( .A(\alu_b[18] ), .Z(\malu/_048_ ) );
BUF_X1 \malu/_517_ ( .A(\malu/_217_ ), .Z(\malu/r[18] ) );
BUF_X1 \malu/_518_ ( .A(\alu_b[19] ), .Z(\malu/_049_ ) );
BUF_X1 \malu/_519_ ( .A(\malu/_218_ ), .Z(\malu/r[19] ) );
BUF_X1 \malu/_520_ ( .A(\alu_b[20] ), .Z(\malu/_051_ ) );
BUF_X1 \malu/_521_ ( .A(\malu/_220_ ), .Z(\malu/r[20] ) );
BUF_X1 \malu/_522_ ( .A(\alu_b[21] ), .Z(\malu/_052_ ) );
BUF_X1 \malu/_523_ ( .A(\malu/_221_ ), .Z(\malu/r[21] ) );
BUF_X1 \malu/_524_ ( .A(\alu_b[22] ), .Z(\malu/_053_ ) );
BUF_X1 \malu/_525_ ( .A(\malu/_222_ ), .Z(\malu/r[22] ) );
BUF_X1 \malu/_526_ ( .A(\alu_b[23] ), .Z(\malu/_054_ ) );
BUF_X1 \malu/_527_ ( .A(\malu/_223_ ), .Z(\malu/r[23] ) );
BUF_X1 \malu/_528_ ( .A(\alu_b[24] ), .Z(\malu/_055_ ) );
BUF_X1 \malu/_529_ ( .A(\malu/_224_ ), .Z(\malu/r[24] ) );
BUF_X1 \malu/_530_ ( .A(\alu_b[25] ), .Z(\malu/_056_ ) );
BUF_X1 \malu/_531_ ( .A(\malu/_225_ ), .Z(\malu/r[25] ) );
BUF_X1 \malu/_532_ ( .A(\alu_b[26] ), .Z(\malu/_057_ ) );
BUF_X1 \malu/_533_ ( .A(\malu/_226_ ), .Z(\malu/r[26] ) );
BUF_X1 \malu/_534_ ( .A(\alu_b[27] ), .Z(\malu/_058_ ) );
BUF_X1 \malu/_535_ ( .A(\malu/_227_ ), .Z(\malu/r[27] ) );
BUF_X1 \malu/_536_ ( .A(\alu_b[28] ), .Z(\malu/_059_ ) );
BUF_X1 \malu/_537_ ( .A(\malu/_228_ ), .Z(\malu/r[28] ) );
BUF_X1 \malu/_538_ ( .A(\alu_b[29] ), .Z(\malu/_060_ ) );
BUF_X1 \malu/_539_ ( .A(\malu/_229_ ), .Z(\malu/r[29] ) );
BUF_X1 \malu/_540_ ( .A(\alu_b[30] ), .Z(\malu/_062_ ) );
BUF_X1 \malu/_541_ ( .A(\malu/_231_ ), .Z(\malu/r[30] ) );
BUF_X1 \malu/_542_ ( .A(\alu_b[31] ), .Z(\malu/_063_ ) );
BUF_X1 \malu/_543_ ( .A(\malu/_232_ ), .Z(\malu/r[31] ) );
BUF_X1 \malu/_544_ ( .A(\alu_ctl[0] ), .Z(\malu/_035_ ) );
BUF_X1 \malu/_545_ ( .A(\alu_ctl[1] ), .Z(\malu/_036_ ) );
BUF_X1 \malu/_546_ ( .A(\alu_ctl[2] ), .Z(\malu/_037_ ) );
BUF_X1 \malu/_547_ ( .A(\alu_ctl[3] ), .Z(\malu/_038_ ) );
BUF_X1 \malu/_548_ ( .A(\malu/_272_ ), .Z(\malu/shift_ctl[0] ) );
BUF_X1 \malu/_549_ ( .A(\malu/_273_ ), .Z(\malu/shift_ctl[1] ) );
BUF_X1 \malu/_550_ ( .A(\malu/_072_ ), .Z(\malu/logic_ctl[0] ) );
BUF_X1 \malu/_551_ ( .A(\malu/_073_ ), .Z(\malu/logic_ctl[1] ) );
BUF_X1 \malu/_552_ ( .A(OF ), .Z(\malu/_001_ ) );
BUF_X1 \malu/_553_ ( .A(\malu/adder_result[31] ), .Z(\malu/_027_ ) );
BUF_X1 \malu/_554_ ( .A(CF ), .Z(\malu/_000_ ) );
BUF_X1 \malu/_555_ ( .A(alu_sign ), .Z(\malu/_306_ ) );
BUF_X1 \malu/_556_ ( .A(\malu/logic_result[0] ), .Z(\malu/_074_ ) );
BUF_X1 \malu/_557_ ( .A(\malu/shift_result[0] ), .Z(\malu/_274_ ) );
BUF_X1 \malu/_558_ ( .A(\malu/adder_result[0] ), .Z(\malu/_003_ ) );
BUF_X1 \malu/_559_ ( .A(\malu/_240_ ), .Z(\alu_result[0] ) );
BUF_X1 \malu/_560_ ( .A(\malu/logic_result[1] ), .Z(\malu/_085_ ) );
BUF_X1 \malu/_561_ ( .A(\malu/shift_result[1] ), .Z(\malu/_285_ ) );
BUF_X1 \malu/_562_ ( .A(\malu/adder_result[1] ), .Z(\malu/_014_ ) );
BUF_X1 \malu/_563_ ( .A(\malu/_251_ ), .Z(\alu_result[1] ) );
BUF_X1 \malu/_564_ ( .A(\malu/logic_result[2] ), .Z(\malu/_096_ ) );
BUF_X1 \malu/_565_ ( .A(\malu/shift_result[2] ), .Z(\malu/_296_ ) );
BUF_X1 \malu/_566_ ( .A(\malu/adder_result[2] ), .Z(\malu/_025_ ) );
BUF_X1 \malu/_567_ ( .A(\malu/_262_ ), .Z(\alu_result[2] ) );
BUF_X1 \malu/_568_ ( .A(\malu/logic_result[3] ), .Z(\malu/_099_ ) );
BUF_X1 \malu/_569_ ( .A(\malu/shift_result[3] ), .Z(\malu/_299_ ) );
BUF_X1 \malu/_570_ ( .A(\malu/adder_result[3] ), .Z(\malu/_028_ ) );
BUF_X1 \malu/_571_ ( .A(\malu/_265_ ), .Z(\alu_result[3] ) );
BUF_X1 \malu/_572_ ( .A(\malu/logic_result[4] ), .Z(\malu/_100_ ) );
BUF_X1 \malu/_573_ ( .A(\malu/shift_result[4] ), .Z(\malu/_300_ ) );
BUF_X1 \malu/_574_ ( .A(\malu/adder_result[4] ), .Z(\malu/_029_ ) );
BUF_X1 \malu/_575_ ( .A(\malu/_266_ ), .Z(\alu_result[4] ) );
BUF_X1 \malu/_576_ ( .A(\malu/logic_result[5] ), .Z(\malu/_101_ ) );
BUF_X1 \malu/_577_ ( .A(\malu/shift_result[5] ), .Z(\malu/_301_ ) );
BUF_X1 \malu/_578_ ( .A(\malu/adder_result[5] ), .Z(\malu/_030_ ) );
BUF_X1 \malu/_579_ ( .A(\malu/_267_ ), .Z(\alu_result[5] ) );
BUF_X1 \malu/_580_ ( .A(\malu/logic_result[6] ), .Z(\malu/_102_ ) );
BUF_X1 \malu/_581_ ( .A(\malu/shift_result[6] ), .Z(\malu/_302_ ) );
BUF_X1 \malu/_582_ ( .A(\malu/adder_result[6] ), .Z(\malu/_031_ ) );
BUF_X1 \malu/_583_ ( .A(\malu/_268_ ), .Z(\alu_result[6] ) );
BUF_X1 \malu/_584_ ( .A(\malu/logic_result[7] ), .Z(\malu/_103_ ) );
BUF_X1 \malu/_585_ ( .A(\malu/shift_result[7] ), .Z(\malu/_303_ ) );
BUF_X1 \malu/_586_ ( .A(\malu/adder_result[7] ), .Z(\malu/_032_ ) );
BUF_X1 \malu/_587_ ( .A(\malu/_269_ ), .Z(\alu_result[7] ) );
BUF_X1 \malu/_588_ ( .A(\malu/logic_result[8] ), .Z(\malu/_104_ ) );
BUF_X1 \malu/_589_ ( .A(\malu/shift_result[8] ), .Z(\malu/_304_ ) );
BUF_X1 \malu/_590_ ( .A(\malu/adder_result[8] ), .Z(\malu/_033_ ) );
BUF_X1 \malu/_591_ ( .A(\malu/_270_ ), .Z(\alu_result[8] ) );
BUF_X1 \malu/_592_ ( .A(\malu/logic_result[9] ), .Z(\malu/_105_ ) );
BUF_X1 \malu/_593_ ( .A(\malu/shift_result[9] ), .Z(\malu/_305_ ) );
BUF_X1 \malu/_594_ ( .A(\malu/adder_result[9] ), .Z(\malu/_034_ ) );
BUF_X1 \malu/_595_ ( .A(\malu/_271_ ), .Z(\alu_result[9] ) );
BUF_X1 \malu/_596_ ( .A(\malu/logic_result[10] ), .Z(\malu/_075_ ) );
BUF_X1 \malu/_597_ ( .A(\malu/shift_result[10] ), .Z(\malu/_275_ ) );
BUF_X1 \malu/_598_ ( .A(\malu/adder_result[10] ), .Z(\malu/_004_ ) );
BUF_X1 \malu/_599_ ( .A(\malu/_241_ ), .Z(\alu_result[10] ) );
BUF_X1 \malu/_600_ ( .A(\malu/logic_result[11] ), .Z(\malu/_076_ ) );
BUF_X1 \malu/_601_ ( .A(\malu/shift_result[11] ), .Z(\malu/_276_ ) );
BUF_X1 \malu/_602_ ( .A(\malu/adder_result[11] ), .Z(\malu/_005_ ) );
BUF_X1 \malu/_603_ ( .A(\malu/_242_ ), .Z(\alu_result[11] ) );
BUF_X1 \malu/_604_ ( .A(\malu/logic_result[12] ), .Z(\malu/_077_ ) );
BUF_X1 \malu/_605_ ( .A(\malu/shift_result[12] ), .Z(\malu/_277_ ) );
BUF_X1 \malu/_606_ ( .A(\malu/adder_result[12] ), .Z(\malu/_006_ ) );
BUF_X1 \malu/_607_ ( .A(\malu/_243_ ), .Z(\alu_result[12] ) );
BUF_X1 \malu/_608_ ( .A(\malu/logic_result[13] ), .Z(\malu/_078_ ) );
BUF_X1 \malu/_609_ ( .A(\malu/shift_result[13] ), .Z(\malu/_278_ ) );
BUF_X1 \malu/_610_ ( .A(\malu/adder_result[13] ), .Z(\malu/_007_ ) );
BUF_X1 \malu/_611_ ( .A(\malu/_244_ ), .Z(\alu_result[13] ) );
BUF_X1 \malu/_612_ ( .A(\malu/logic_result[14] ), .Z(\malu/_079_ ) );
BUF_X1 \malu/_613_ ( .A(\malu/shift_result[14] ), .Z(\malu/_279_ ) );
BUF_X1 \malu/_614_ ( .A(\malu/adder_result[14] ), .Z(\malu/_008_ ) );
BUF_X1 \malu/_615_ ( .A(\malu/_245_ ), .Z(\alu_result[14] ) );
BUF_X1 \malu/_616_ ( .A(\malu/logic_result[15] ), .Z(\malu/_080_ ) );
BUF_X1 \malu/_617_ ( .A(\malu/shift_result[15] ), .Z(\malu/_280_ ) );
BUF_X1 \malu/_618_ ( .A(\malu/adder_result[15] ), .Z(\malu/_009_ ) );
BUF_X1 \malu/_619_ ( .A(\malu/_246_ ), .Z(\alu_result[15] ) );
BUF_X1 \malu/_620_ ( .A(\malu/logic_result[16] ), .Z(\malu/_081_ ) );
BUF_X1 \malu/_621_ ( .A(\malu/shift_result[16] ), .Z(\malu/_281_ ) );
BUF_X1 \malu/_622_ ( .A(\malu/adder_result[16] ), .Z(\malu/_010_ ) );
BUF_X1 \malu/_623_ ( .A(\malu/_247_ ), .Z(\alu_result[16] ) );
BUF_X1 \malu/_624_ ( .A(\malu/logic_result[17] ), .Z(\malu/_082_ ) );
BUF_X1 \malu/_625_ ( .A(\malu/shift_result[17] ), .Z(\malu/_282_ ) );
BUF_X1 \malu/_626_ ( .A(\malu/adder_result[17] ), .Z(\malu/_011_ ) );
BUF_X1 \malu/_627_ ( .A(\malu/_248_ ), .Z(\alu_result[17] ) );
BUF_X1 \malu/_628_ ( .A(\malu/logic_result[18] ), .Z(\malu/_083_ ) );
BUF_X1 \malu/_629_ ( .A(\malu/shift_result[18] ), .Z(\malu/_283_ ) );
BUF_X1 \malu/_630_ ( .A(\malu/adder_result[18] ), .Z(\malu/_012_ ) );
BUF_X1 \malu/_631_ ( .A(\malu/_249_ ), .Z(\alu_result[18] ) );
BUF_X1 \malu/_632_ ( .A(\malu/logic_result[19] ), .Z(\malu/_084_ ) );
BUF_X1 \malu/_633_ ( .A(\malu/shift_result[19] ), .Z(\malu/_284_ ) );
BUF_X1 \malu/_634_ ( .A(\malu/adder_result[19] ), .Z(\malu/_013_ ) );
BUF_X1 \malu/_635_ ( .A(\malu/_250_ ), .Z(\alu_result[19] ) );
BUF_X1 \malu/_636_ ( .A(\malu/logic_result[20] ), .Z(\malu/_086_ ) );
BUF_X1 \malu/_637_ ( .A(\malu/shift_result[20] ), .Z(\malu/_286_ ) );
BUF_X1 \malu/_638_ ( .A(\malu/adder_result[20] ), .Z(\malu/_015_ ) );
BUF_X1 \malu/_639_ ( .A(\malu/_252_ ), .Z(\alu_result[20] ) );
BUF_X1 \malu/_640_ ( .A(\malu/logic_result[21] ), .Z(\malu/_087_ ) );
BUF_X1 \malu/_641_ ( .A(\malu/shift_result[21] ), .Z(\malu/_287_ ) );
BUF_X1 \malu/_642_ ( .A(\malu/adder_result[21] ), .Z(\malu/_016_ ) );
BUF_X1 \malu/_643_ ( .A(\malu/_253_ ), .Z(\alu_result[21] ) );
BUF_X1 \malu/_644_ ( .A(\malu/logic_result[22] ), .Z(\malu/_088_ ) );
BUF_X1 \malu/_645_ ( .A(\malu/shift_result[22] ), .Z(\malu/_288_ ) );
BUF_X1 \malu/_646_ ( .A(\malu/adder_result[22] ), .Z(\malu/_017_ ) );
BUF_X1 \malu/_647_ ( .A(\malu/_254_ ), .Z(\alu_result[22] ) );
BUF_X1 \malu/_648_ ( .A(\malu/logic_result[23] ), .Z(\malu/_089_ ) );
BUF_X1 \malu/_649_ ( .A(\malu/shift_result[23] ), .Z(\malu/_289_ ) );
BUF_X1 \malu/_650_ ( .A(\malu/adder_result[23] ), .Z(\malu/_018_ ) );
BUF_X1 \malu/_651_ ( .A(\malu/_255_ ), .Z(\alu_result[23] ) );
BUF_X1 \malu/_652_ ( .A(\malu/logic_result[24] ), .Z(\malu/_090_ ) );
BUF_X1 \malu/_653_ ( .A(\malu/shift_result[24] ), .Z(\malu/_290_ ) );
BUF_X1 \malu/_654_ ( .A(\malu/adder_result[24] ), .Z(\malu/_019_ ) );
BUF_X1 \malu/_655_ ( .A(\malu/_256_ ), .Z(\alu_result[24] ) );
BUF_X1 \malu/_656_ ( .A(\malu/logic_result[25] ), .Z(\malu/_091_ ) );
BUF_X1 \malu/_657_ ( .A(\malu/shift_result[25] ), .Z(\malu/_291_ ) );
BUF_X1 \malu/_658_ ( .A(\malu/adder_result[25] ), .Z(\malu/_020_ ) );
BUF_X1 \malu/_659_ ( .A(\malu/_257_ ), .Z(\alu_result[25] ) );
BUF_X1 \malu/_660_ ( .A(\malu/logic_result[26] ), .Z(\malu/_092_ ) );
BUF_X1 \malu/_661_ ( .A(\malu/shift_result[26] ), .Z(\malu/_292_ ) );
BUF_X1 \malu/_662_ ( .A(\malu/adder_result[26] ), .Z(\malu/_021_ ) );
BUF_X1 \malu/_663_ ( .A(\malu/_258_ ), .Z(\alu_result[26] ) );
BUF_X1 \malu/_664_ ( .A(\malu/logic_result[27] ), .Z(\malu/_093_ ) );
BUF_X1 \malu/_665_ ( .A(\malu/shift_result[27] ), .Z(\malu/_293_ ) );
BUF_X1 \malu/_666_ ( .A(\malu/adder_result[27] ), .Z(\malu/_022_ ) );
BUF_X1 \malu/_667_ ( .A(\malu/_259_ ), .Z(\alu_result[27] ) );
BUF_X1 \malu/_668_ ( .A(\malu/logic_result[28] ), .Z(\malu/_094_ ) );
BUF_X1 \malu/_669_ ( .A(\malu/shift_result[28] ), .Z(\malu/_294_ ) );
BUF_X1 \malu/_670_ ( .A(\malu/adder_result[28] ), .Z(\malu/_023_ ) );
BUF_X1 \malu/_671_ ( .A(\malu/_260_ ), .Z(\alu_result[28] ) );
BUF_X1 \malu/_672_ ( .A(\malu/logic_result[29] ), .Z(\malu/_095_ ) );
BUF_X1 \malu/_673_ ( .A(\malu/shift_result[29] ), .Z(\malu/_295_ ) );
BUF_X1 \malu/_674_ ( .A(\malu/adder_result[29] ), .Z(\malu/_024_ ) );
BUF_X1 \malu/_675_ ( .A(\malu/_261_ ), .Z(\alu_result[29] ) );
BUF_X1 \malu/_676_ ( .A(\malu/logic_result[30] ), .Z(\malu/_097_ ) );
BUF_X1 \malu/_677_ ( .A(\malu/shift_result[30] ), .Z(\malu/_297_ ) );
BUF_X1 \malu/_678_ ( .A(\malu/adder_result[30] ), .Z(\malu/_026_ ) );
BUF_X1 \malu/_679_ ( .A(\malu/_263_ ), .Z(\alu_result[30] ) );
BUF_X1 \malu/_680_ ( .A(\malu/logic_result[31] ), .Z(\malu/_098_ ) );
BUF_X1 \malu/_681_ ( .A(\malu/shift_result[31] ), .Z(\malu/_298_ ) );
BUF_X1 \malu/_682_ ( .A(\malu/_264_ ), .Z(\alu_result[31] ) );
BUF_X1 \malu/_683_ ( .A(ZF ), .Z(\malu/_002_ ) );
BUF_X1 \malu/_684_ ( .A(\malu/_071_ ), .Z(branch ) );
XOR2_X2 \malu/Adder/_324_ ( .A(\malu/Adder/_032_ ), .B(\malu/Adder/_000_ ), .Z(\malu/Adder/_066_ ) );
XOR2_X1 \malu/Adder/_325_ ( .A(\malu/Adder/_066_ ), .B(\malu/Adder/_064_ ), .Z(\malu/Adder/_291_ ) );
AND2_X4 \malu/Adder/_326_ ( .A1(\malu/Adder/_066_ ), .A2(\malu/Adder/_064_ ), .ZN(\malu/Adder/_067_ ) );
AND2_X1 \malu/Adder/_327_ ( .A1(\malu/Adder/_032_ ), .A2(\malu/Adder/_000_ ), .ZN(\malu/Adder/_068_ ) );
NOR2_X4 \malu/Adder/_328_ ( .A1(\malu/Adder/_067_ ), .A2(\malu/Adder/_068_ ), .ZN(\malu/Adder/_069_ ) );
XOR2_X1 \malu/Adder/_329_ ( .A(\malu/Adder/_043_ ), .B(\malu/Adder/_011_ ), .Z(\malu/Adder/_070_ ) );
XNOR2_X1 \malu/Adder/_330_ ( .A(\malu/Adder/_069_ ), .B(\malu/Adder/_070_ ), .ZN(\malu/Adder/_302_ ) );
AND2_X1 \malu/Adder/_331_ ( .A1(\malu/Adder/_043_ ), .A2(\malu/Adder/_011_ ), .ZN(\malu/Adder/_071_ ) );
NOR2_X1 \malu/Adder/_332_ ( .A1(\malu/Adder/_043_ ), .A2(\malu/Adder/_011_ ), .ZN(\malu/Adder/_072_ ) );
NOR3_X4 \malu/Adder/_333_ ( .A1(\malu/Adder/_069_ ), .A2(\malu/Adder/_071_ ), .A3(\malu/Adder/_072_ ), .ZN(\malu/Adder/_073_ ) );
XOR2_X1 \malu/Adder/_334_ ( .A(\malu/Adder/_054_ ), .B(\malu/Adder/_022_ ), .Z(\malu/Adder/_074_ ) );
OR3_X1 \malu/Adder/_335_ ( .A1(\malu/Adder/_073_ ), .A2(\malu/Adder/_071_ ), .A3(\malu/Adder/_074_ ), .ZN(\malu/Adder/_075_ ) );
OAI21_X1 \malu/Adder/_336_ ( .A(\malu/Adder/_074_ ), .B1(\malu/Adder/_073_ ), .B2(\malu/Adder/_071_ ), .ZN(\malu/Adder/_076_ ) );
AND2_X1 \malu/Adder/_337_ ( .A1(\malu/Adder/_075_ ), .A2(\malu/Adder/_076_ ), .ZN(\malu/Adder/_313_ ) );
AND2_X1 \malu/Adder/_338_ ( .A1(\malu/Adder/_054_ ), .A2(\malu/Adder/_022_ ), .ZN(\malu/Adder/_077_ ) );
INV_X1 \malu/Adder/_339_ ( .A(\malu/Adder/_077_ ), .ZN(\malu/Adder/_078_ ) );
NAND2_X1 \malu/Adder/_340_ ( .A1(\malu/Adder/_076_ ), .A2(\malu/Adder/_078_ ), .ZN(\malu/Adder/_079_ ) );
XOR2_X1 \malu/Adder/_341_ ( .A(\malu/Adder/_057_ ), .B(\malu/Adder/_025_ ), .Z(\malu/Adder/_080_ ) );
XNOR2_X1 \malu/Adder/_342_ ( .A(\malu/Adder/_079_ ), .B(\malu/Adder/_080_ ), .ZN(\malu/Adder/_081_ ) );
INV_X1 \malu/Adder/_343_ ( .A(\malu/Adder/_081_ ), .ZN(\malu/Adder/_316_ ) );
OAI211_X2 \malu/Adder/_344_ ( .A(\malu/Adder/_074_ ), .B(\malu/Adder/_080_ ), .C1(\malu/Adder/_073_ ), .C2(\malu/Adder/_071_ ), .ZN(\malu/Adder/_082_ ) );
AND2_X1 \malu/Adder/_345_ ( .A1(\malu/Adder/_080_ ), .A2(\malu/Adder/_077_ ), .ZN(\malu/Adder/_083_ ) );
AOI21_X1 \malu/Adder/_346_ ( .A(\malu/Adder/_083_ ), .B1(\malu/Adder/_057_ ), .B2(\malu/Adder/_025_ ), .ZN(\malu/Adder/_084_ ) );
AND2_X4 \malu/Adder/_347_ ( .A1(\malu/Adder/_082_ ), .A2(\malu/Adder/_084_ ), .ZN(\malu/Adder/_085_ ) );
XOR2_X1 \malu/Adder/_348_ ( .A(\malu/Adder/_058_ ), .B(\malu/Adder/_026_ ), .Z(\malu/Adder/_086_ ) );
XNOR2_X1 \malu/Adder/_349_ ( .A(\malu/Adder/_085_ ), .B(\malu/Adder/_086_ ), .ZN(\malu/Adder/_317_ ) );
NOR2_X1 \malu/Adder/_350_ ( .A1(\malu/Adder/_058_ ), .A2(\malu/Adder/_026_ ), .ZN(\malu/Adder/_087_ ) );
AND2_X1 \malu/Adder/_351_ ( .A1(\malu/Adder/_058_ ), .A2(\malu/Adder/_026_ ), .ZN(\malu/Adder/_088_ ) );
NOR3_X1 \malu/Adder/_352_ ( .A1(\malu/Adder/_085_ ), .A2(\malu/Adder/_087_ ), .A3(\malu/Adder/_088_ ), .ZN(\malu/Adder/_089_ ) );
OR2_X1 \malu/Adder/_353_ ( .A1(\malu/Adder/_089_ ), .A2(\malu/Adder/_088_ ), .ZN(\malu/Adder/_090_ ) );
XOR2_X2 \malu/Adder/_354_ ( .A(\malu/Adder/_059_ ), .B(\malu/Adder/_027_ ), .Z(\malu/Adder/_091_ ) );
XNOR2_X1 \malu/Adder/_355_ ( .A(\malu/Adder/_090_ ), .B(\malu/Adder/_091_ ), .ZN(\malu/Adder/_092_ ) );
INV_X1 \malu/Adder/_356_ ( .A(\malu/Adder/_092_ ), .ZN(\malu/Adder/_318_ ) );
INV_X4 \malu/Adder/_357_ ( .A(\malu/Adder/_085_ ), .ZN(\malu/Adder/_093_ ) );
AND2_X1 \malu/Adder/_358_ ( .A1(\malu/Adder/_086_ ), .A2(\malu/Adder/_091_ ), .ZN(\malu/Adder/_094_ ) );
NAND2_X1 \malu/Adder/_359_ ( .A1(\malu/Adder/_093_ ), .A2(\malu/Adder/_094_ ), .ZN(\malu/Adder/_095_ ) );
AND2_X4 \malu/Adder/_360_ ( .A1(\malu/Adder/_091_ ), .A2(\malu/Adder/_088_ ), .ZN(\malu/Adder/_096_ ) );
AOI21_X4 \malu/Adder/_361_ ( .A(\malu/Adder/_096_ ), .B1(\malu/Adder/_059_ ), .B2(\malu/Adder/_027_ ), .ZN(\malu/Adder/_097_ ) );
NAND2_X1 \malu/Adder/_362_ ( .A1(\malu/Adder/_095_ ), .A2(\malu/Adder/_097_ ), .ZN(\malu/Adder/_098_ ) );
XOR2_X1 \malu/Adder/_363_ ( .A(\malu/Adder/_060_ ), .B(\malu/Adder/_028_ ), .Z(\malu/Adder/_099_ ) );
INV_X1 \malu/Adder/_364_ ( .A(\malu/Adder/_099_ ), .ZN(\malu/Adder/_100_ ) );
XNOR2_X1 \malu/Adder/_365_ ( .A(\malu/Adder/_098_ ), .B(\malu/Adder/_100_ ), .ZN(\malu/Adder/_319_ ) );
NAND2_X1 \malu/Adder/_366_ ( .A1(\malu/Adder/_098_ ), .A2(\malu/Adder/_099_ ), .ZN(\malu/Adder/_101_ ) );
NAND2_X1 \malu/Adder/_367_ ( .A1(\malu/Adder/_060_ ), .A2(\malu/Adder/_028_ ), .ZN(\malu/Adder/_102_ ) );
NAND2_X1 \malu/Adder/_368_ ( .A1(\malu/Adder/_101_ ), .A2(\malu/Adder/_102_ ), .ZN(\malu/Adder/_103_ ) );
XOR2_X1 \malu/Adder/_369_ ( .A(\malu/Adder/_061_ ), .B(\malu/Adder/_029_ ), .Z(\malu/Adder/_104_ ) );
INV_X1 \malu/Adder/_370_ ( .A(\malu/Adder/_104_ ), .ZN(\malu/Adder/_105_ ) );
XNOR2_X1 \malu/Adder/_371_ ( .A(\malu/Adder/_103_ ), .B(\malu/Adder/_105_ ), .ZN(\malu/Adder/_320_ ) );
NAND4_X4 \malu/Adder/_372_ ( .A1(\malu/Adder/_093_ ), .A2(\malu/Adder/_094_ ), .A3(\malu/Adder/_099_ ), .A4(\malu/Adder/_104_ ), .ZN(\malu/Adder/_106_ ) );
AND3_X1 \malu/Adder/_373_ ( .A1(\malu/Adder/_104_ ), .A2(\malu/Adder/_060_ ), .A3(\malu/Adder/_028_ ), .ZN(\malu/Adder/_107_ ) );
NOR3_X1 \malu/Adder/_374_ ( .A1(\malu/Adder/_097_ ), .A2(\malu/Adder/_100_ ), .A3(\malu/Adder/_105_ ), .ZN(\malu/Adder/_108_ ) );
AOI211_X2 \malu/Adder/_375_ ( .A(\malu/Adder/_107_ ), .B(\malu/Adder/_108_ ), .C1(\malu/Adder/_061_ ), .C2(\malu/Adder/_029_ ), .ZN(\malu/Adder/_109_ ) );
AND2_X2 \malu/Adder/_376_ ( .A1(\malu/Adder/_106_ ), .A2(\malu/Adder/_109_ ), .ZN(\malu/Adder/_110_ ) );
XOR2_X1 \malu/Adder/_377_ ( .A(\malu/Adder/_062_ ), .B(\malu/Adder/_030_ ), .Z(\malu/Adder/_111_ ) );
XNOR2_X1 \malu/Adder/_378_ ( .A(\malu/Adder/_110_ ), .B(\malu/Adder/_111_ ), .ZN(\malu/Adder/_321_ ) );
NOR2_X1 \malu/Adder/_379_ ( .A1(\malu/Adder/_062_ ), .A2(\malu/Adder/_030_ ), .ZN(\malu/Adder/_112_ ) );
AND2_X1 \malu/Adder/_380_ ( .A1(\malu/Adder/_062_ ), .A2(\malu/Adder/_030_ ), .ZN(\malu/Adder/_113_ ) );
NOR3_X1 \malu/Adder/_381_ ( .A1(\malu/Adder/_110_ ), .A2(\malu/Adder/_112_ ), .A3(\malu/Adder/_113_ ), .ZN(\malu/Adder/_114_ ) );
NOR2_X1 \malu/Adder/_382_ ( .A1(\malu/Adder/_114_ ), .A2(\malu/Adder/_113_ ), .ZN(\malu/Adder/_115_ ) );
XOR2_X2 \malu/Adder/_383_ ( .A(\malu/Adder/_063_ ), .B(\malu/Adder/_031_ ), .Z(\malu/Adder/_116_ ) );
XNOR2_X1 \malu/Adder/_384_ ( .A(\malu/Adder/_115_ ), .B(\malu/Adder/_116_ ), .ZN(\malu/Adder/_322_ ) );
NAND2_X1 \malu/Adder/_385_ ( .A1(\malu/Adder/_111_ ), .A2(\malu/Adder/_116_ ), .ZN(\malu/Adder/_117_ ) );
OR2_X1 \malu/Adder/_386_ ( .A1(\malu/Adder/_110_ ), .A2(\malu/Adder/_117_ ), .ZN(\malu/Adder/_118_ ) );
AND2_X2 \malu/Adder/_387_ ( .A1(\malu/Adder/_116_ ), .A2(\malu/Adder/_113_ ), .ZN(\malu/Adder/_119_ ) );
AOI21_X2 \malu/Adder/_388_ ( .A(\malu/Adder/_119_ ), .B1(\malu/Adder/_063_ ), .B2(\malu/Adder/_031_ ), .ZN(\malu/Adder/_120_ ) );
NAND2_X1 \malu/Adder/_389_ ( .A1(\malu/Adder/_118_ ), .A2(\malu/Adder/_120_ ), .ZN(\malu/Adder/_121_ ) );
XOR2_X1 \malu/Adder/_390_ ( .A(\malu/Adder/_033_ ), .B(\malu/Adder/_001_ ), .Z(\malu/Adder/_122_ ) );
INV_X1 \malu/Adder/_391_ ( .A(\malu/Adder/_122_ ), .ZN(\malu/Adder/_123_ ) );
XNOR2_X1 \malu/Adder/_392_ ( .A(\malu/Adder/_121_ ), .B(\malu/Adder/_123_ ), .ZN(\malu/Adder/_292_ ) );
NAND2_X1 \malu/Adder/_393_ ( .A1(\malu/Adder/_121_ ), .A2(\malu/Adder/_122_ ), .ZN(\malu/Adder/_124_ ) );
NAND2_X1 \malu/Adder/_394_ ( .A1(\malu/Adder/_033_ ), .A2(\malu/Adder/_001_ ), .ZN(\malu/Adder/_125_ ) );
NAND2_X1 \malu/Adder/_395_ ( .A1(\malu/Adder/_124_ ), .A2(\malu/Adder/_125_ ), .ZN(\malu/Adder/_126_ ) );
XOR2_X1 \malu/Adder/_396_ ( .A(\malu/Adder/_034_ ), .B(\malu/Adder/_002_ ), .Z(\malu/Adder/_127_ ) );
XNOR2_X1 \malu/Adder/_397_ ( .A(\malu/Adder/_126_ ), .B(\malu/Adder/_127_ ), .ZN(\malu/Adder/_128_ ) );
INV_X1 \malu/Adder/_398_ ( .A(\malu/Adder/_128_ ), .ZN(\malu/Adder/_293_ ) );
AND2_X1 \malu/Adder/_399_ ( .A1(\malu/Adder/_111_ ), .A2(\malu/Adder/_116_ ), .ZN(\malu/Adder/_129_ ) );
AND3_X1 \malu/Adder/_400_ ( .A1(\malu/Adder/_129_ ), .A2(\malu/Adder/_122_ ), .A3(\malu/Adder/_127_ ), .ZN(\malu/Adder/_130_ ) );
INV_X1 \malu/Adder/_401_ ( .A(\malu/Adder/_130_ ), .ZN(\malu/Adder/_131_ ) );
OR2_X4 \malu/Adder/_402_ ( .A1(\malu/Adder/_110_ ), .A2(\malu/Adder/_131_ ), .ZN(\malu/Adder/_132_ ) );
NOR2_X1 \malu/Adder/_403_ ( .A1(\malu/Adder/_034_ ), .A2(\malu/Adder/_002_ ), .ZN(\malu/Adder/_133_ ) );
AND2_X1 \malu/Adder/_404_ ( .A1(\malu/Adder/_034_ ), .A2(\malu/Adder/_002_ ), .ZN(\malu/Adder/_134_ ) );
NOR4_X2 \malu/Adder/_405_ ( .A1(\malu/Adder/_123_ ), .A2(\malu/Adder/_120_ ), .A3(\malu/Adder/_133_ ), .A4(\malu/Adder/_134_ ), .ZN(\malu/Adder/_135_ ) );
NOR3_X1 \malu/Adder/_406_ ( .A1(\malu/Adder/_134_ ), .A2(\malu/Adder/_133_ ), .A3(\malu/Adder/_125_ ), .ZN(\malu/Adder/_136_ ) );
NOR3_X2 \malu/Adder/_407_ ( .A1(\malu/Adder/_135_ ), .A2(\malu/Adder/_134_ ), .A3(\malu/Adder/_136_ ), .ZN(\malu/Adder/_137_ ) );
AND2_X4 \malu/Adder/_408_ ( .A1(\malu/Adder/_132_ ), .A2(\malu/Adder/_137_ ), .ZN(\malu/Adder/_138_ ) );
XOR2_X1 \malu/Adder/_409_ ( .A(\malu/Adder/_035_ ), .B(\malu/Adder/_003_ ), .Z(\malu/Adder/_139_ ) );
XNOR2_X1 \malu/Adder/_410_ ( .A(\malu/Adder/_138_ ), .B(\malu/Adder/_139_ ), .ZN(\malu/Adder/_294_ ) );
INV_X1 \malu/Adder/_411_ ( .A(\malu/Adder/_139_ ), .ZN(\malu/Adder/_140_ ) );
OR2_X1 \malu/Adder/_412_ ( .A1(\malu/Adder/_138_ ), .A2(\malu/Adder/_140_ ), .ZN(\malu/Adder/_141_ ) );
NAND2_X1 \malu/Adder/_413_ ( .A1(\malu/Adder/_035_ ), .A2(\malu/Adder/_003_ ), .ZN(\malu/Adder/_142_ ) );
NAND2_X1 \malu/Adder/_414_ ( .A1(\malu/Adder/_141_ ), .A2(\malu/Adder/_142_ ), .ZN(\malu/Adder/_143_ ) );
AND2_X1 \malu/Adder/_415_ ( .A1(\malu/Adder/_036_ ), .A2(\malu/Adder/_004_ ), .ZN(\malu/Adder/_144_ ) );
NOR2_X4 \malu/Adder/_416_ ( .A1(\malu/Adder/_036_ ), .A2(\malu/Adder/_004_ ), .ZN(\malu/Adder/_145_ ) );
NOR2_X1 \malu/Adder/_417_ ( .A1(\malu/Adder/_144_ ), .A2(\malu/Adder/_145_ ), .ZN(\malu/Adder/_146_ ) );
XNOR2_X1 \malu/Adder/_418_ ( .A(\malu/Adder/_143_ ), .B(\malu/Adder/_146_ ), .ZN(\malu/Adder/_147_ ) );
INV_X1 \malu/Adder/_419_ ( .A(\malu/Adder/_147_ ), .ZN(\malu/Adder/_295_ ) );
NOR4_X4 \malu/Adder/_420_ ( .A1(\malu/Adder/_138_ ), .A2(\malu/Adder/_140_ ), .A3(\malu/Adder/_144_ ), .A4(\malu/Adder/_145_ ), .ZN(\malu/Adder/_148_ ) );
NOR3_X1 \malu/Adder/_421_ ( .A1(\malu/Adder/_144_ ), .A2(\malu/Adder/_145_ ), .A3(\malu/Adder/_142_ ), .ZN(\malu/Adder/_149_ ) );
OR2_X1 \malu/Adder/_422_ ( .A1(\malu/Adder/_149_ ), .A2(\malu/Adder/_144_ ), .ZN(\malu/Adder/_150_ ) );
NOR2_X4 \malu/Adder/_423_ ( .A1(\malu/Adder/_148_ ), .A2(\malu/Adder/_150_ ), .ZN(\malu/Adder/_151_ ) );
XOR2_X1 \malu/Adder/_424_ ( .A(\malu/Adder/_037_ ), .B(\malu/Adder/_005_ ), .Z(\malu/Adder/_152_ ) );
XNOR2_X1 \malu/Adder/_425_ ( .A(\malu/Adder/_151_ ), .B(\malu/Adder/_152_ ), .ZN(\malu/Adder/_296_ ) );
NOR2_X1 \malu/Adder/_426_ ( .A1(\malu/Adder/_037_ ), .A2(\malu/Adder/_005_ ), .ZN(\malu/Adder/_153_ ) );
AND2_X1 \malu/Adder/_427_ ( .A1(\malu/Adder/_037_ ), .A2(\malu/Adder/_005_ ), .ZN(\malu/Adder/_154_ ) );
NOR3_X2 \malu/Adder/_428_ ( .A1(\malu/Adder/_151_ ), .A2(\malu/Adder/_153_ ), .A3(\malu/Adder/_154_ ), .ZN(\malu/Adder/_155_ ) );
NOR2_X1 \malu/Adder/_429_ ( .A1(\malu/Adder/_155_ ), .A2(\malu/Adder/_154_ ), .ZN(\malu/Adder/_156_ ) );
XOR2_X1 \malu/Adder/_430_ ( .A(\malu/Adder/_038_ ), .B(\malu/Adder/_006_ ), .Z(\malu/Adder/_157_ ) );
XNOR2_X1 \malu/Adder/_431_ ( .A(\malu/Adder/_156_ ), .B(\malu/Adder/_157_ ), .ZN(\malu/Adder/_297_ ) );
AND2_X1 \malu/Adder/_432_ ( .A1(\malu/Adder/_152_ ), .A2(\malu/Adder/_157_ ), .ZN(\malu/Adder/_158_ ) );
AND3_X1 \malu/Adder/_433_ ( .A1(\malu/Adder/_158_ ), .A2(\malu/Adder/_139_ ), .A3(\malu/Adder/_146_ ), .ZN(\malu/Adder/_159_ ) );
INV_X1 \malu/Adder/_434_ ( .A(\malu/Adder/_159_ ), .ZN(\malu/Adder/_160_ ) );
AOI211_X4 \malu/Adder/_435_ ( .A(\malu/Adder/_131_ ), .B(\malu/Adder/_160_ ), .C1(\malu/Adder/_106_ ), .C2(\malu/Adder/_109_ ), .ZN(\malu/Adder/_161_ ) );
NOR2_X2 \malu/Adder/_436_ ( .A1(\malu/Adder/_137_ ), .A2(\malu/Adder/_160_ ), .ZN(\malu/Adder/_162_ ) );
AND2_X1 \malu/Adder/_437_ ( .A1(\malu/Adder/_038_ ), .A2(\malu/Adder/_006_ ), .ZN(\malu/Adder/_163_ ) );
AND2_X1 \malu/Adder/_438_ ( .A1(\malu/Adder/_150_ ), .A2(\malu/Adder/_158_ ), .ZN(\malu/Adder/_164_ ) );
AND2_X1 \malu/Adder/_439_ ( .A1(\malu/Adder/_157_ ), .A2(\malu/Adder/_154_ ), .ZN(\malu/Adder/_165_ ) );
NOR4_X4 \malu/Adder/_440_ ( .A1(\malu/Adder/_162_ ), .A2(\malu/Adder/_163_ ), .A3(\malu/Adder/_164_ ), .A4(\malu/Adder/_165_ ), .ZN(\malu/Adder/_166_ ) );
INV_X2 \malu/Adder/_441_ ( .A(\malu/Adder/_166_ ), .ZN(\malu/Adder/_167_ ) );
XOR2_X1 \malu/Adder/_442_ ( .A(\malu/Adder/_039_ ), .B(\malu/Adder/_007_ ), .Z(\malu/Adder/_168_ ) );
OR3_X4 \malu/Adder/_443_ ( .A1(\malu/Adder/_161_ ), .A2(\malu/Adder/_167_ ), .A3(\malu/Adder/_168_ ), .ZN(\malu/Adder/_169_ ) );
OAI21_X1 \malu/Adder/_444_ ( .A(\malu/Adder/_168_ ), .B1(\malu/Adder/_161_ ), .B2(\malu/Adder/_167_ ), .ZN(\malu/Adder/_170_ ) );
AND2_X4 \malu/Adder/_445_ ( .A1(\malu/Adder/_169_ ), .A2(\malu/Adder/_170_ ), .ZN(\malu/Adder/_298_ ) );
AND2_X1 \malu/Adder/_446_ ( .A1(\malu/Adder/_039_ ), .A2(\malu/Adder/_007_ ), .ZN(\malu/Adder/_171_ ) );
INV_X1 \malu/Adder/_447_ ( .A(\malu/Adder/_171_ ), .ZN(\malu/Adder/_172_ ) );
NAND2_X1 \malu/Adder/_448_ ( .A1(\malu/Adder/_170_ ), .A2(\malu/Adder/_172_ ), .ZN(\malu/Adder/_173_ ) );
XOR2_X1 \malu/Adder/_449_ ( .A(\malu/Adder/_040_ ), .B(\malu/Adder/_008_ ), .Z(\malu/Adder/_174_ ) );
XNOR2_X1 \malu/Adder/_450_ ( .A(\malu/Adder/_173_ ), .B(\malu/Adder/_174_ ), .ZN(\malu/Adder/_175_ ) );
INV_X1 \malu/Adder/_451_ ( .A(\malu/Adder/_175_ ), .ZN(\malu/Adder/_299_ ) );
AND2_X1 \malu/Adder/_452_ ( .A1(\malu/Adder/_168_ ), .A2(\malu/Adder/_174_ ), .ZN(\malu/Adder/_176_ ) );
OAI21_X1 \malu/Adder/_453_ ( .A(\malu/Adder/_176_ ), .B1(\malu/Adder/_161_ ), .B2(\malu/Adder/_167_ ), .ZN(\malu/Adder/_177_ ) );
AND2_X1 \malu/Adder/_454_ ( .A1(\malu/Adder/_174_ ), .A2(\malu/Adder/_171_ ), .ZN(\malu/Adder/_178_ ) );
AOI21_X1 \malu/Adder/_455_ ( .A(\malu/Adder/_178_ ), .B1(\malu/Adder/_040_ ), .B2(\malu/Adder/_008_ ), .ZN(\malu/Adder/_179_ ) );
NAND2_X1 \malu/Adder/_456_ ( .A1(\malu/Adder/_177_ ), .A2(\malu/Adder/_179_ ), .ZN(\malu/Adder/_180_ ) );
XOR2_X1 \malu/Adder/_457_ ( .A(\malu/Adder/_041_ ), .B(\malu/Adder/_009_ ), .Z(\malu/Adder/_181_ ) );
XOR2_X1 \malu/Adder/_458_ ( .A(\malu/Adder/_180_ ), .B(\malu/Adder/_181_ ), .Z(\malu/Adder/_300_ ) );
NAND2_X1 \malu/Adder/_459_ ( .A1(\malu/Adder/_180_ ), .A2(\malu/Adder/_181_ ), .ZN(\malu/Adder/_182_ ) );
AND2_X1 \malu/Adder/_460_ ( .A1(\malu/Adder/_041_ ), .A2(\malu/Adder/_009_ ), .ZN(\malu/Adder/_183_ ) );
INV_X1 \malu/Adder/_461_ ( .A(\malu/Adder/_183_ ), .ZN(\malu/Adder/_184_ ) );
AND2_X1 \malu/Adder/_462_ ( .A1(\malu/Adder/_182_ ), .A2(\malu/Adder/_184_ ), .ZN(\malu/Adder/_185_ ) );
XOR2_X1 \malu/Adder/_463_ ( .A(\malu/Adder/_042_ ), .B(\malu/Adder/_010_ ), .Z(\malu/Adder/_186_ ) );
XNOR2_X1 \malu/Adder/_464_ ( .A(\malu/Adder/_185_ ), .B(\malu/Adder/_186_ ), .ZN(\malu/Adder/_301_ ) );
XOR2_X1 \malu/Adder/_465_ ( .A(\malu/Adder/_044_ ), .B(\malu/Adder/_012_ ), .Z(\malu/Adder/_187_ ) );
AND2_X1 \malu/Adder/_466_ ( .A1(\malu/Adder/_181_ ), .A2(\malu/Adder/_186_ ), .ZN(\malu/Adder/_188_ ) );
AND2_X1 \malu/Adder/_467_ ( .A1(\malu/Adder/_188_ ), .A2(\malu/Adder/_176_ ), .ZN(\malu/Adder/_189_ ) );
INV_X1 \malu/Adder/_468_ ( .A(\malu/Adder/_189_ ), .ZN(\malu/Adder/_190_ ) );
INV_X2 \malu/Adder/_469_ ( .A(\malu/Adder/_161_ ), .ZN(\malu/Adder/_191_ ) );
AOI21_X2 \malu/Adder/_470_ ( .A(\malu/Adder/_190_ ), .B1(\malu/Adder/_191_ ), .B2(\malu/Adder/_166_ ), .ZN(\malu/Adder/_192_ ) );
AND2_X1 \malu/Adder/_471_ ( .A1(\malu/Adder/_186_ ), .A2(\malu/Adder/_183_ ), .ZN(\malu/Adder/_193_ ) );
AOI21_X1 \malu/Adder/_472_ ( .A(\malu/Adder/_193_ ), .B1(\malu/Adder/_042_ ), .B2(\malu/Adder/_010_ ), .ZN(\malu/Adder/_194_ ) );
INV_X1 \malu/Adder/_473_ ( .A(\malu/Adder/_188_ ), .ZN(\malu/Adder/_195_ ) );
OAI21_X1 \malu/Adder/_474_ ( .A(\malu/Adder/_194_ ), .B1(\malu/Adder/_179_ ), .B2(\malu/Adder/_195_ ), .ZN(\malu/Adder/_196_ ) );
OAI21_X1 \malu/Adder/_475_ ( .A(\malu/Adder/_187_ ), .B1(\malu/Adder/_192_ ), .B2(\malu/Adder/_196_ ), .ZN(\malu/Adder/_197_ ) );
OR3_X1 \malu/Adder/_476_ ( .A1(\malu/Adder/_192_ ), .A2(\malu/Adder/_196_ ), .A3(\malu/Adder/_187_ ), .ZN(\malu/Adder/_198_ ) );
AND2_X2 \malu/Adder/_477_ ( .A1(\malu/Adder/_197_ ), .A2(\malu/Adder/_198_ ), .ZN(\malu/Adder/_303_ ) );
NAND2_X1 \malu/Adder/_478_ ( .A1(\malu/Adder/_044_ ), .A2(\malu/Adder/_012_ ), .ZN(\malu/Adder/_199_ ) );
AND2_X1 \malu/Adder/_479_ ( .A1(\malu/Adder/_197_ ), .A2(\malu/Adder/_199_ ), .ZN(\malu/Adder/_200_ ) );
AND2_X1 \malu/Adder/_480_ ( .A1(\malu/Adder/_045_ ), .A2(\malu/Adder/_013_ ), .ZN(\malu/Adder/_201_ ) );
NOR2_X1 \malu/Adder/_481_ ( .A1(\malu/Adder/_045_ ), .A2(\malu/Adder/_013_ ), .ZN(\malu/Adder/_202_ ) );
NOR2_X1 \malu/Adder/_482_ ( .A1(\malu/Adder/_201_ ), .A2(\malu/Adder/_202_ ), .ZN(\malu/Adder/_203_ ) );
XNOR2_X1 \malu/Adder/_483_ ( .A(\malu/Adder/_200_ ), .B(\malu/Adder/_203_ ), .ZN(\malu/Adder/_304_ ) );
AND2_X1 \malu/Adder/_484_ ( .A1(\malu/Adder/_187_ ), .A2(\malu/Adder/_203_ ), .ZN(\malu/Adder/_204_ ) );
OAI21_X1 \malu/Adder/_485_ ( .A(\malu/Adder/_204_ ), .B1(\malu/Adder/_192_ ), .B2(\malu/Adder/_196_ ), .ZN(\malu/Adder/_205_ ) );
NOR3_X1 \malu/Adder/_486_ ( .A1(\malu/Adder/_201_ ), .A2(\malu/Adder/_202_ ), .A3(\malu/Adder/_199_ ), .ZN(\malu/Adder/_206_ ) );
NOR2_X1 \malu/Adder/_487_ ( .A1(\malu/Adder/_206_ ), .A2(\malu/Adder/_201_ ), .ZN(\malu/Adder/_207_ ) );
AND2_X1 \malu/Adder/_488_ ( .A1(\malu/Adder/_205_ ), .A2(\malu/Adder/_207_ ), .ZN(\malu/Adder/_208_ ) );
XOR2_X1 \malu/Adder/_489_ ( .A(\malu/Adder/_046_ ), .B(\malu/Adder/_014_ ), .Z(\malu/Adder/_209_ ) );
XNOR2_X1 \malu/Adder/_490_ ( .A(\malu/Adder/_208_ ), .B(\malu/Adder/_209_ ), .ZN(\malu/Adder/_305_ ) );
NOR2_X1 \malu/Adder/_491_ ( .A1(\malu/Adder/_046_ ), .A2(\malu/Adder/_014_ ), .ZN(\malu/Adder/_210_ ) );
AND2_X1 \malu/Adder/_492_ ( .A1(\malu/Adder/_046_ ), .A2(\malu/Adder/_014_ ), .ZN(\malu/Adder/_211_ ) );
NOR3_X1 \malu/Adder/_493_ ( .A1(\malu/Adder/_208_ ), .A2(\malu/Adder/_210_ ), .A3(\malu/Adder/_211_ ), .ZN(\malu/Adder/_212_ ) );
NOR2_X1 \malu/Adder/_494_ ( .A1(\malu/Adder/_212_ ), .A2(\malu/Adder/_211_ ), .ZN(\malu/Adder/_213_ ) );
XOR2_X1 \malu/Adder/_495_ ( .A(\malu/Adder/_047_ ), .B(\malu/Adder/_015_ ), .Z(\malu/Adder/_214_ ) );
XNOR2_X1 \malu/Adder/_496_ ( .A(\malu/Adder/_213_ ), .B(\malu/Adder/_214_ ), .ZN(\malu/Adder/_306_ ) );
AND2_X1 \malu/Adder/_497_ ( .A1(\malu/Adder/_209_ ), .A2(\malu/Adder/_214_ ), .ZN(\malu/Adder/_215_ ) );
AND2_X1 \malu/Adder/_498_ ( .A1(\malu/Adder/_215_ ), .A2(\malu/Adder/_204_ ), .ZN(\malu/Adder/_216_ ) );
OAI211_X2 \malu/Adder/_499_ ( .A(\malu/Adder/_189_ ), .B(\malu/Adder/_216_ ), .C1(\malu/Adder/_161_ ), .C2(\malu/Adder/_167_ ), .ZN(\malu/Adder/_217_ ) );
NAND2_X1 \malu/Adder/_500_ ( .A1(\malu/Adder/_196_ ), .A2(\malu/Adder/_216_ ), .ZN(\malu/Adder/_218_ ) );
OAI21_X1 \malu/Adder/_501_ ( .A(\malu/Adder/_215_ ), .B1(\malu/Adder/_201_ ), .B2(\malu/Adder/_206_ ), .ZN(\malu/Adder/_219_ ) );
AND2_X1 \malu/Adder/_502_ ( .A1(\malu/Adder/_214_ ), .A2(\malu/Adder/_211_ ), .ZN(\malu/Adder/_220_ ) );
AOI21_X1 \malu/Adder/_503_ ( .A(\malu/Adder/_220_ ), .B1(\malu/Adder/_047_ ), .B2(\malu/Adder/_015_ ), .ZN(\malu/Adder/_221_ ) );
AND3_X1 \malu/Adder/_504_ ( .A1(\malu/Adder/_218_ ), .A2(\malu/Adder/_219_ ), .A3(\malu/Adder/_221_ ), .ZN(\malu/Adder/_222_ ) );
AND2_X4 \malu/Adder/_505_ ( .A1(\malu/Adder/_217_ ), .A2(\malu/Adder/_222_ ), .ZN(\malu/Adder/_223_ ) );
XOR2_X1 \malu/Adder/_506_ ( .A(\malu/Adder/_048_ ), .B(\malu/Adder/_016_ ), .Z(\malu/Adder/_224_ ) );
XNOR2_X2 \malu/Adder/_507_ ( .A(\malu/Adder/_223_ ), .B(\malu/Adder/_224_ ), .ZN(\malu/Adder/_307_ ) );
INV_X1 \malu/Adder/_508_ ( .A(\malu/Adder/_224_ ), .ZN(\malu/Adder/_225_ ) );
OR2_X1 \malu/Adder/_509_ ( .A1(\malu/Adder/_223_ ), .A2(\malu/Adder/_225_ ), .ZN(\malu/Adder/_226_ ) );
NAND2_X1 \malu/Adder/_510_ ( .A1(\malu/Adder/_048_ ), .A2(\malu/Adder/_016_ ), .ZN(\malu/Adder/_227_ ) );
AND2_X1 \malu/Adder/_511_ ( .A1(\malu/Adder/_226_ ), .A2(\malu/Adder/_227_ ), .ZN(\malu/Adder/_228_ ) );
AND2_X1 \malu/Adder/_512_ ( .A1(\malu/Adder/_049_ ), .A2(\malu/Adder/_017_ ), .ZN(\malu/Adder/_229_ ) );
NOR2_X1 \malu/Adder/_513_ ( .A1(\malu/Adder/_049_ ), .A2(\malu/Adder/_017_ ), .ZN(\malu/Adder/_230_ ) );
NOR2_X1 \malu/Adder/_514_ ( .A1(\malu/Adder/_229_ ), .A2(\malu/Adder/_230_ ), .ZN(\malu/Adder/_231_ ) );
XNOR2_X1 \malu/Adder/_515_ ( .A(\malu/Adder/_228_ ), .B(\malu/Adder/_231_ ), .ZN(\malu/Adder/_308_ ) );
NOR4_X1 \malu/Adder/_516_ ( .A1(\malu/Adder/_223_ ), .A2(\malu/Adder/_225_ ), .A3(\malu/Adder/_230_ ), .A4(\malu/Adder/_229_ ), .ZN(\malu/Adder/_232_ ) );
NOR3_X1 \malu/Adder/_517_ ( .A1(\malu/Adder/_229_ ), .A2(\malu/Adder/_230_ ), .A3(\malu/Adder/_227_ ), .ZN(\malu/Adder/_233_ ) );
OR2_X1 \malu/Adder/_518_ ( .A1(\malu/Adder/_233_ ), .A2(\malu/Adder/_229_ ), .ZN(\malu/Adder/_234_ ) );
NOR2_X1 \malu/Adder/_519_ ( .A1(\malu/Adder/_232_ ), .A2(\malu/Adder/_234_ ), .ZN(\malu/Adder/_235_ ) );
XOR2_X1 \malu/Adder/_520_ ( .A(\malu/Adder/_050_ ), .B(\malu/Adder/_018_ ), .Z(\malu/Adder/_236_ ) );
XNOR2_X1 \malu/Adder/_521_ ( .A(\malu/Adder/_235_ ), .B(\malu/Adder/_236_ ), .ZN(\malu/Adder/_309_ ) );
OAI21_X1 \malu/Adder/_522_ ( .A(\malu/Adder/_236_ ), .B1(\malu/Adder/_232_ ), .B2(\malu/Adder/_234_ ), .ZN(\malu/Adder/_237_ ) );
AND2_X1 \malu/Adder/_523_ ( .A1(\malu/Adder/_050_ ), .A2(\malu/Adder/_018_ ), .ZN(\malu/Adder/_238_ ) );
INV_X1 \malu/Adder/_524_ ( .A(\malu/Adder/_238_ ), .ZN(\malu/Adder/_239_ ) );
NAND2_X1 \malu/Adder/_525_ ( .A1(\malu/Adder/_237_ ), .A2(\malu/Adder/_239_ ), .ZN(\malu/Adder/_240_ ) );
XOR2_X1 \malu/Adder/_526_ ( .A(\malu/Adder/_051_ ), .B(\malu/Adder/_019_ ), .Z(\malu/Adder/_241_ ) );
XNOR2_X1 \malu/Adder/_527_ ( .A(\malu/Adder/_240_ ), .B(\malu/Adder/_241_ ), .ZN(\malu/Adder/_242_ ) );
INV_X1 \malu/Adder/_528_ ( .A(\malu/Adder/_242_ ), .ZN(\malu/Adder/_310_ ) );
AND2_X1 \malu/Adder/_529_ ( .A1(\malu/Adder/_236_ ), .A2(\malu/Adder/_241_ ), .ZN(\malu/Adder/_243_ ) );
NAND3_X1 \malu/Adder/_530_ ( .A1(\malu/Adder/_243_ ), .A2(\malu/Adder/_224_ ), .A3(\malu/Adder/_231_ ), .ZN(\malu/Adder/_244_ ) );
OR2_X1 \malu/Adder/_531_ ( .A1(\malu/Adder/_223_ ), .A2(\malu/Adder/_244_ ), .ZN(\malu/Adder/_245_ ) );
AND2_X1 \malu/Adder/_532_ ( .A1(\malu/Adder/_234_ ), .A2(\malu/Adder/_243_ ), .ZN(\malu/Adder/_246_ ) );
AND2_X1 \malu/Adder/_533_ ( .A1(\malu/Adder/_051_ ), .A2(\malu/Adder/_019_ ), .ZN(\malu/Adder/_247_ ) );
AND2_X1 \malu/Adder/_534_ ( .A1(\malu/Adder/_241_ ), .A2(\malu/Adder/_238_ ), .ZN(\malu/Adder/_248_ ) );
NOR3_X1 \malu/Adder/_535_ ( .A1(\malu/Adder/_246_ ), .A2(\malu/Adder/_247_ ), .A3(\malu/Adder/_248_ ), .ZN(\malu/Adder/_249_ ) );
NAND2_X1 \malu/Adder/_536_ ( .A1(\malu/Adder/_245_ ), .A2(\malu/Adder/_249_ ), .ZN(\malu/Adder/_250_ ) );
XOR2_X1 \malu/Adder/_537_ ( .A(\malu/Adder/_052_ ), .B(\malu/Adder/_020_ ), .Z(\malu/Adder/_251_ ) );
XOR2_X1 \malu/Adder/_538_ ( .A(\malu/Adder/_250_ ), .B(\malu/Adder/_251_ ), .Z(\malu/Adder/_311_ ) );
NAND2_X1 \malu/Adder/_539_ ( .A1(\malu/Adder/_250_ ), .A2(\malu/Adder/_251_ ), .ZN(\malu/Adder/_252_ ) );
AND2_X1 \malu/Adder/_540_ ( .A1(\malu/Adder/_052_ ), .A2(\malu/Adder/_020_ ), .ZN(\malu/Adder/_253_ ) );
INV_X1 \malu/Adder/_541_ ( .A(\malu/Adder/_253_ ), .ZN(\malu/Adder/_254_ ) );
NAND2_X1 \malu/Adder/_542_ ( .A1(\malu/Adder/_252_ ), .A2(\malu/Adder/_254_ ), .ZN(\malu/Adder/_255_ ) );
XOR2_X1 \malu/Adder/_543_ ( .A(\malu/Adder/_053_ ), .B(\malu/Adder/_021_ ), .Z(\malu/Adder/_256_ ) );
XNOR2_X1 \malu/Adder/_544_ ( .A(\malu/Adder/_255_ ), .B(\malu/Adder/_256_ ), .ZN(\malu/Adder/_257_ ) );
INV_X1 \malu/Adder/_545_ ( .A(\malu/Adder/_257_ ), .ZN(\malu/Adder/_312_ ) );
AND2_X1 \malu/Adder/_546_ ( .A1(\malu/Adder/_251_ ), .A2(\malu/Adder/_256_ ), .ZN(\malu/Adder/_258_ ) );
NAND2_X1 \malu/Adder/_547_ ( .A1(\malu/Adder/_250_ ), .A2(\malu/Adder/_258_ ), .ZN(\malu/Adder/_259_ ) );
AND2_X1 \malu/Adder/_548_ ( .A1(\malu/Adder/_256_ ), .A2(\malu/Adder/_253_ ), .ZN(\malu/Adder/_260_ ) );
AOI21_X1 \malu/Adder/_549_ ( .A(\malu/Adder/_260_ ), .B1(\malu/Adder/_053_ ), .B2(\malu/Adder/_021_ ), .ZN(\malu/Adder/_261_ ) );
XOR2_X1 \malu/Adder/_550_ ( .A(\malu/Adder/_055_ ), .B(\malu/Adder/_023_ ), .Z(\malu/Adder/_262_ ) );
INV_X1 \malu/Adder/_551_ ( .A(\malu/Adder/_262_ ), .ZN(\malu/Adder/_263_ ) );
AND3_X1 \malu/Adder/_552_ ( .A1(\malu/Adder/_259_ ), .A2(\malu/Adder/_261_ ), .A3(\malu/Adder/_263_ ), .ZN(\malu/Adder/_264_ ) );
AOI21_X1 \malu/Adder/_553_ ( .A(\malu/Adder/_263_ ), .B1(\malu/Adder/_259_ ), .B2(\malu/Adder/_261_ ), .ZN(\malu/Adder/_265_ ) );
NOR2_X1 \malu/Adder/_554_ ( .A1(\malu/Adder/_264_ ), .A2(\malu/Adder/_265_ ), .ZN(\malu/Adder/_314_ ) );
AND2_X1 \malu/Adder/_555_ ( .A1(\malu/Adder/_055_ ), .A2(\malu/Adder/_023_ ), .ZN(\malu/Adder/_266_ ) );
NOR2_X1 \malu/Adder/_556_ ( .A1(\malu/Adder/_265_ ), .A2(\malu/Adder/_266_ ), .ZN(\malu/Adder/_267_ ) );
AND2_X1 \malu/Adder/_557_ ( .A1(\malu/Adder/_056_ ), .A2(\malu/Adder/_024_ ), .ZN(\malu/Adder/_268_ ) );
NOR2_X1 \malu/Adder/_558_ ( .A1(\malu/Adder/_056_ ), .A2(\malu/Adder/_024_ ), .ZN(\malu/Adder/_269_ ) );
NOR2_X1 \malu/Adder/_559_ ( .A1(\malu/Adder/_268_ ), .A2(\malu/Adder/_269_ ), .ZN(\malu/Adder/_270_ ) );
XNOR2_X1 \malu/Adder/_560_ ( .A(\malu/Adder/_267_ ), .B(\malu/Adder/_270_ ), .ZN(\malu/Adder/_315_ ) );
XNOR2_X1 \malu/Adder/_561_ ( .A(\malu/Adder/_267_ ), .B(\malu/Adder/_024_ ), .ZN(\malu/Adder/_271_ ) );
INV_X1 \malu/Adder/_562_ ( .A(\malu/Adder/_270_ ), .ZN(\malu/Adder/_272_ ) );
AND2_X1 \malu/Adder/_563_ ( .A1(\malu/Adder/_271_ ), .A2(\malu/Adder/_272_ ), .ZN(\malu/Adder/_290_ ) );
OR4_X2 \malu/Adder/_564_ ( .A1(\malu/Adder/_297_ ), .A2(\malu/Adder/_300_ ), .A3(\malu/Adder/_303_ ), .A4(\malu/Adder/_307_ ), .ZN(\malu/Adder/_273_ ) );
NOR3_X2 \malu/Adder/_565_ ( .A1(\malu/Adder/_273_ ), .A2(\malu/Adder/_301_ ), .A3(\malu/Adder/_304_ ), .ZN(\malu/Adder/_274_ ) );
NOR4_X4 \malu/Adder/_566_ ( .A1(\malu/Adder/_294_ ), .A2(\malu/Adder/_322_ ), .A3(\malu/Adder/_292_ ), .A4(\malu/Adder/_298_ ), .ZN(\malu/Adder/_275_ ) );
NOR4_X1 \malu/Adder/_567_ ( .A1(\malu/Adder/_317_ ), .A2(\malu/Adder/_291_ ), .A3(\malu/Adder/_302_ ), .A4(\malu/Adder/_313_ ), .ZN(\malu/Adder/_276_ ) );
NAND3_X1 \malu/Adder/_568_ ( .A1(\malu/Adder/_092_ ), .A2(\malu/Adder/_081_ ), .A3(\malu/Adder/_276_ ), .ZN(\malu/Adder/_277_ ) );
NOR4_X1 \malu/Adder/_569_ ( .A1(\malu/Adder/_320_ ), .A2(\malu/Adder/_277_ ), .A3(\malu/Adder/_319_ ), .A4(\malu/Adder/_321_ ), .ZN(\malu/Adder/_278_ ) );
NAND2_X1 \malu/Adder/_570_ ( .A1(\malu/Adder/_275_ ), .A2(\malu/Adder/_278_ ), .ZN(\malu/Adder/_279_ ) );
NOR3_X1 \malu/Adder/_571_ ( .A1(\malu/Adder/_279_ ), .A2(\malu/Adder/_296_ ), .A3(\malu/Adder/_293_ ), .ZN(\malu/Adder/_280_ ) );
AND3_X1 \malu/Adder/_572_ ( .A1(\malu/Adder/_280_ ), .A2(\malu/Adder/_147_ ), .A3(\malu/Adder/_175_ ), .ZN(\malu/Adder/_281_ ) );
NAND2_X1 \malu/Adder/_573_ ( .A1(\malu/Adder/_274_ ), .A2(\malu/Adder/_281_ ), .ZN(\malu/Adder/_282_ ) );
OR4_X2 \malu/Adder/_574_ ( .A1(\malu/Adder/_305_ ), .A2(\malu/Adder/_282_ ), .A3(\malu/Adder/_309_ ), .A4(\malu/Adder/_311_ ), .ZN(\malu/Adder/_283_ ) );
OR4_X2 \malu/Adder/_575_ ( .A1(\malu/Adder/_310_ ), .A2(\malu/Adder/_283_ ), .A3(\malu/Adder/_312_ ), .A4(\malu/Adder/_314_ ), .ZN(\malu/Adder/_284_ ) );
NOR4_X1 \malu/Adder/_576_ ( .A1(\malu/Adder/_284_ ), .A2(\malu/Adder/_306_ ), .A3(\malu/Adder/_308_ ), .A4(\malu/Adder/_315_ ), .ZN(\malu/Adder/_323_ ) );
NAND3_X1 \malu/Adder/_577_ ( .A1(\malu/Adder/_258_ ), .A2(\malu/Adder/_262_ ), .A3(\malu/Adder/_270_ ), .ZN(\malu/Adder/_285_ ) );
OR3_X1 \malu/Adder/_578_ ( .A1(\malu/Adder/_223_ ), .A2(\malu/Adder/_244_ ), .A3(\malu/Adder/_285_ ), .ZN(\malu/Adder/_286_ ) );
OR2_X1 \malu/Adder/_579_ ( .A1(\malu/Adder/_249_ ), .A2(\malu/Adder/_285_ ), .ZN(\malu/Adder/_287_ ) );
OR3_X1 \malu/Adder/_580_ ( .A1(\malu/Adder/_261_ ), .A2(\malu/Adder/_263_ ), .A3(\malu/Adder/_272_ ), .ZN(\malu/Adder/_288_ ) );
AOI21_X1 \malu/Adder/_581_ ( .A(\malu/Adder/_268_ ), .B1(\malu/Adder/_270_ ), .B2(\malu/Adder/_266_ ), .ZN(\malu/Adder/_289_ ) );
NAND4_X1 \malu/Adder/_582_ ( .A1(\malu/Adder/_286_ ), .A2(\malu/Adder/_287_ ), .A3(\malu/Adder/_288_ ), .A4(\malu/Adder/_289_ ), .ZN(\malu/Adder/_065_ ) );
BUF_X1 \malu/Adder/_583_ ( .A(\malu/r[0] ), .Z(\malu/Adder/_032_ ) );
BUF_X1 \malu/Adder/_584_ ( .A(\alu_a[0] ), .Z(\malu/Adder/_000_ ) );
BUF_X1 \malu/Adder/_585_ ( .A(alu_sub ), .Z(\malu/Adder/_064_ ) );
BUF_X1 \malu/Adder/_586_ ( .A(\malu/Adder/_291_ ), .Z(\malu/adder_result[0] ) );
BUF_X1 \malu/Adder/_587_ ( .A(\malu/r[1] ), .Z(\malu/Adder/_043_ ) );
BUF_X1 \malu/Adder/_588_ ( .A(\alu_a[1] ), .Z(\malu/Adder/_011_ ) );
BUF_X1 \malu/Adder/_589_ ( .A(\malu/Adder/_302_ ), .Z(\malu/adder_result[1] ) );
BUF_X1 \malu/Adder/_590_ ( .A(\malu/r[2] ), .Z(\malu/Adder/_054_ ) );
BUF_X1 \malu/Adder/_591_ ( .A(\alu_a[2] ), .Z(\malu/Adder/_022_ ) );
BUF_X1 \malu/Adder/_592_ ( .A(\malu/Adder/_313_ ), .Z(\malu/adder_result[2] ) );
BUF_X1 \malu/Adder/_593_ ( .A(\malu/r[3] ), .Z(\malu/Adder/_057_ ) );
BUF_X1 \malu/Adder/_594_ ( .A(\alu_a[3] ), .Z(\malu/Adder/_025_ ) );
BUF_X1 \malu/Adder/_595_ ( .A(\malu/Adder/_316_ ), .Z(\malu/adder_result[3] ) );
BUF_X1 \malu/Adder/_596_ ( .A(\malu/r[4] ), .Z(\malu/Adder/_058_ ) );
BUF_X1 \malu/Adder/_597_ ( .A(\alu_a[4] ), .Z(\malu/Adder/_026_ ) );
BUF_X1 \malu/Adder/_598_ ( .A(\malu/Adder/_317_ ), .Z(\malu/adder_result[4] ) );
BUF_X1 \malu/Adder/_599_ ( .A(\malu/r[5] ), .Z(\malu/Adder/_059_ ) );
BUF_X1 \malu/Adder/_600_ ( .A(\alu_a[5] ), .Z(\malu/Adder/_027_ ) );
BUF_X1 \malu/Adder/_601_ ( .A(\malu/Adder/_318_ ), .Z(\malu/adder_result[5] ) );
BUF_X1 \malu/Adder/_602_ ( .A(\malu/r[6] ), .Z(\malu/Adder/_060_ ) );
BUF_X1 \malu/Adder/_603_ ( .A(\alu_a[6] ), .Z(\malu/Adder/_028_ ) );
BUF_X1 \malu/Adder/_604_ ( .A(\malu/Adder/_319_ ), .Z(\malu/adder_result[6] ) );
BUF_X1 \malu/Adder/_605_ ( .A(\malu/r[7] ), .Z(\malu/Adder/_061_ ) );
BUF_X1 \malu/Adder/_606_ ( .A(\alu_a[7] ), .Z(\malu/Adder/_029_ ) );
BUF_X1 \malu/Adder/_607_ ( .A(\malu/Adder/_320_ ), .Z(\malu/adder_result[7] ) );
BUF_X1 \malu/Adder/_608_ ( .A(\malu/r[8] ), .Z(\malu/Adder/_062_ ) );
BUF_X1 \malu/Adder/_609_ ( .A(\alu_a[8] ), .Z(\malu/Adder/_030_ ) );
BUF_X1 \malu/Adder/_610_ ( .A(\malu/Adder/_321_ ), .Z(\malu/adder_result[8] ) );
BUF_X1 \malu/Adder/_611_ ( .A(\malu/r[9] ), .Z(\malu/Adder/_063_ ) );
BUF_X1 \malu/Adder/_612_ ( .A(\alu_a[9] ), .Z(\malu/Adder/_031_ ) );
BUF_X1 \malu/Adder/_613_ ( .A(\malu/Adder/_322_ ), .Z(\malu/adder_result[9] ) );
BUF_X1 \malu/Adder/_614_ ( .A(\malu/r[10] ), .Z(\malu/Adder/_033_ ) );
BUF_X1 \malu/Adder/_615_ ( .A(\alu_a[10] ), .Z(\malu/Adder/_001_ ) );
BUF_X1 \malu/Adder/_616_ ( .A(\malu/Adder/_292_ ), .Z(\malu/adder_result[10] ) );
BUF_X1 \malu/Adder/_617_ ( .A(\malu/r[11] ), .Z(\malu/Adder/_034_ ) );
BUF_X1 \malu/Adder/_618_ ( .A(\alu_a[11] ), .Z(\malu/Adder/_002_ ) );
BUF_X1 \malu/Adder/_619_ ( .A(\malu/Adder/_293_ ), .Z(\malu/adder_result[11] ) );
BUF_X1 \malu/Adder/_620_ ( .A(\malu/r[12] ), .Z(\malu/Adder/_035_ ) );
BUF_X1 \malu/Adder/_621_ ( .A(\alu_a[12] ), .Z(\malu/Adder/_003_ ) );
BUF_X1 \malu/Adder/_622_ ( .A(\malu/Adder/_294_ ), .Z(\malu/adder_result[12] ) );
BUF_X1 \malu/Adder/_623_ ( .A(\malu/r[13] ), .Z(\malu/Adder/_036_ ) );
BUF_X1 \malu/Adder/_624_ ( .A(\alu_a[13] ), .Z(\malu/Adder/_004_ ) );
BUF_X1 \malu/Adder/_625_ ( .A(\malu/Adder/_295_ ), .Z(\malu/adder_result[13] ) );
BUF_X1 \malu/Adder/_626_ ( .A(\malu/r[14] ), .Z(\malu/Adder/_037_ ) );
BUF_X1 \malu/Adder/_627_ ( .A(\alu_a[14] ), .Z(\malu/Adder/_005_ ) );
BUF_X1 \malu/Adder/_628_ ( .A(\malu/Adder/_296_ ), .Z(\malu/adder_result[14] ) );
BUF_X1 \malu/Adder/_629_ ( .A(\malu/r[15] ), .Z(\malu/Adder/_038_ ) );
BUF_X1 \malu/Adder/_630_ ( .A(\alu_a[15] ), .Z(\malu/Adder/_006_ ) );
BUF_X1 \malu/Adder/_631_ ( .A(\malu/Adder/_297_ ), .Z(\malu/adder_result[15] ) );
BUF_X1 \malu/Adder/_632_ ( .A(\malu/r[16] ), .Z(\malu/Adder/_039_ ) );
BUF_X1 \malu/Adder/_633_ ( .A(\alu_a[16] ), .Z(\malu/Adder/_007_ ) );
BUF_X1 \malu/Adder/_634_ ( .A(\malu/Adder/_298_ ), .Z(\malu/adder_result[16] ) );
BUF_X1 \malu/Adder/_635_ ( .A(\malu/r[17] ), .Z(\malu/Adder/_040_ ) );
BUF_X1 \malu/Adder/_636_ ( .A(\alu_a[17] ), .Z(\malu/Adder/_008_ ) );
BUF_X1 \malu/Adder/_637_ ( .A(\malu/Adder/_299_ ), .Z(\malu/adder_result[17] ) );
BUF_X1 \malu/Adder/_638_ ( .A(\malu/r[18] ), .Z(\malu/Adder/_041_ ) );
BUF_X1 \malu/Adder/_639_ ( .A(\alu_a[18] ), .Z(\malu/Adder/_009_ ) );
BUF_X1 \malu/Adder/_640_ ( .A(\malu/Adder/_300_ ), .Z(\malu/adder_result[18] ) );
BUF_X1 \malu/Adder/_641_ ( .A(\malu/r[19] ), .Z(\malu/Adder/_042_ ) );
BUF_X1 \malu/Adder/_642_ ( .A(\alu_a[19] ), .Z(\malu/Adder/_010_ ) );
BUF_X1 \malu/Adder/_643_ ( .A(\malu/Adder/_301_ ), .Z(\malu/adder_result[19] ) );
BUF_X1 \malu/Adder/_644_ ( .A(\malu/r[20] ), .Z(\malu/Adder/_044_ ) );
BUF_X1 \malu/Adder/_645_ ( .A(\alu_a[20] ), .Z(\malu/Adder/_012_ ) );
BUF_X1 \malu/Adder/_646_ ( .A(\malu/Adder/_303_ ), .Z(\malu/adder_result[20] ) );
BUF_X1 \malu/Adder/_647_ ( .A(\malu/r[21] ), .Z(\malu/Adder/_045_ ) );
BUF_X1 \malu/Adder/_648_ ( .A(\alu_a[21] ), .Z(\malu/Adder/_013_ ) );
BUF_X1 \malu/Adder/_649_ ( .A(\malu/Adder/_304_ ), .Z(\malu/adder_result[21] ) );
BUF_X1 \malu/Adder/_650_ ( .A(\malu/r[22] ), .Z(\malu/Adder/_046_ ) );
BUF_X1 \malu/Adder/_651_ ( .A(\alu_a[22] ), .Z(\malu/Adder/_014_ ) );
BUF_X1 \malu/Adder/_652_ ( .A(\malu/Adder/_305_ ), .Z(\malu/adder_result[22] ) );
BUF_X1 \malu/Adder/_653_ ( .A(\malu/r[23] ), .Z(\malu/Adder/_047_ ) );
BUF_X1 \malu/Adder/_654_ ( .A(\alu_a[23] ), .Z(\malu/Adder/_015_ ) );
BUF_X1 \malu/Adder/_655_ ( .A(\malu/Adder/_306_ ), .Z(\malu/adder_result[23] ) );
BUF_X1 \malu/Adder/_656_ ( .A(\malu/r[24] ), .Z(\malu/Adder/_048_ ) );
BUF_X1 \malu/Adder/_657_ ( .A(\alu_a[24] ), .Z(\malu/Adder/_016_ ) );
BUF_X1 \malu/Adder/_658_ ( .A(\malu/Adder/_307_ ), .Z(\malu/adder_result[24] ) );
BUF_X1 \malu/Adder/_659_ ( .A(\malu/r[25] ), .Z(\malu/Adder/_049_ ) );
BUF_X1 \malu/Adder/_660_ ( .A(\alu_a[25] ), .Z(\malu/Adder/_017_ ) );
BUF_X1 \malu/Adder/_661_ ( .A(\malu/Adder/_308_ ), .Z(\malu/adder_result[25] ) );
BUF_X1 \malu/Adder/_662_ ( .A(\malu/r[26] ), .Z(\malu/Adder/_050_ ) );
BUF_X1 \malu/Adder/_663_ ( .A(\alu_a[26] ), .Z(\malu/Adder/_018_ ) );
BUF_X1 \malu/Adder/_664_ ( .A(\malu/Adder/_309_ ), .Z(\malu/adder_result[26] ) );
BUF_X1 \malu/Adder/_665_ ( .A(\malu/r[27] ), .Z(\malu/Adder/_051_ ) );
BUF_X1 \malu/Adder/_666_ ( .A(\alu_a[27] ), .Z(\malu/Adder/_019_ ) );
BUF_X1 \malu/Adder/_667_ ( .A(\malu/Adder/_310_ ), .Z(\malu/adder_result[27] ) );
BUF_X1 \malu/Adder/_668_ ( .A(\malu/r[28] ), .Z(\malu/Adder/_052_ ) );
BUF_X1 \malu/Adder/_669_ ( .A(\alu_a[28] ), .Z(\malu/Adder/_020_ ) );
BUF_X1 \malu/Adder/_670_ ( .A(\malu/Adder/_311_ ), .Z(\malu/adder_result[28] ) );
BUF_X1 \malu/Adder/_671_ ( .A(\malu/r[29] ), .Z(\malu/Adder/_053_ ) );
BUF_X1 \malu/Adder/_672_ ( .A(\alu_a[29] ), .Z(\malu/Adder/_021_ ) );
BUF_X1 \malu/Adder/_673_ ( .A(\malu/Adder/_312_ ), .Z(\malu/adder_result[29] ) );
BUF_X1 \malu/Adder/_674_ ( .A(\malu/r[30] ), .Z(\malu/Adder/_055_ ) );
BUF_X1 \malu/Adder/_675_ ( .A(\alu_a[30] ), .Z(\malu/Adder/_023_ ) );
BUF_X1 \malu/Adder/_676_ ( .A(\malu/Adder/_314_ ), .Z(\malu/adder_result[30] ) );
BUF_X1 \malu/Adder/_677_ ( .A(\malu/r[31] ), .Z(\malu/Adder/_056_ ) );
BUF_X1 \malu/Adder/_678_ ( .A(\alu_a[31] ), .Z(\malu/Adder/_024_ ) );
BUF_X1 \malu/Adder/_679_ ( .A(\malu/Adder/_315_ ), .Z(\malu/adder_result[31] ) );
BUF_X1 \malu/Adder/_680_ ( .A(\malu/Adder/_290_ ), .Z(OF ) );
BUF_X1 \malu/Adder/_681_ ( .A(\malu/Adder/_323_ ), .Z(ZF ) );
BUF_X1 \malu/Adder/_682_ ( .A(\malu/Adder/_065_ ), .Z(CF ) );
NAND2_X1 \malu/Logic/_202_ ( .A1(\malu/Logic/_032_ ), .A2(\malu/Logic/_000_ ), .ZN(\malu/Logic/_201_ ) );
AOI21_X1 \malu/Logic/_203_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_201_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_098_ ) );
NAND2_X4 \malu/Logic/_204_ ( .A1(\malu/Logic/_064_ ), .A2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_099_ ) );
BUF_X4 \malu/Logic/_205_ ( .A(\malu/Logic/_099_ ), .Z(\malu/Logic/_100_ ) );
AOI21_X2 \malu/Logic/_206_ ( .A(\malu/Logic/_000_ ), .B1(\malu/Logic/_100_ ), .B2(\malu/Logic/_032_ ), .ZN(\malu/Logic/_101_ ) );
OR2_X4 \malu/Logic/_207_ ( .A1(\malu/Logic/_064_ ), .A2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_102_ ) );
OAI22_X1 \malu/Logic/_208_ ( .A1(\malu/Logic/_098_ ), .A2(\malu/Logic/_101_ ), .B1(\malu/Logic/_201_ ), .B2(\malu/Logic/_102_ ), .ZN(\malu/Logic/_066_ ) );
NAND2_X1 \malu/Logic/_209_ ( .A1(\malu/Logic/_043_ ), .A2(\malu/Logic/_011_ ), .ZN(\malu/Logic/_103_ ) );
AOI21_X1 \malu/Logic/_210_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_103_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_104_ ) );
AOI21_X1 \malu/Logic/_211_ ( .A(\malu/Logic/_011_ ), .B1(\malu/Logic/_100_ ), .B2(\malu/Logic/_043_ ), .ZN(\malu/Logic/_105_ ) );
BUF_X4 \malu/Logic/_212_ ( .A(\malu/Logic/_102_ ), .Z(\malu/Logic/_106_ ) );
OAI22_X1 \malu/Logic/_213_ ( .A1(\malu/Logic/_104_ ), .A2(\malu/Logic/_105_ ), .B1(\malu/Logic/_106_ ), .B2(\malu/Logic/_103_ ), .ZN(\malu/Logic/_077_ ) );
NAND2_X1 \malu/Logic/_214_ ( .A1(\malu/Logic/_054_ ), .A2(\malu/Logic/_022_ ), .ZN(\malu/Logic/_107_ ) );
AOI21_X1 \malu/Logic/_215_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_107_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_108_ ) );
AOI21_X1 \malu/Logic/_216_ ( .A(\malu/Logic/_022_ ), .B1(\malu/Logic/_100_ ), .B2(\malu/Logic/_054_ ), .ZN(\malu/Logic/_109_ ) );
OAI22_X1 \malu/Logic/_217_ ( .A1(\malu/Logic/_108_ ), .A2(\malu/Logic/_109_ ), .B1(\malu/Logic/_106_ ), .B2(\malu/Logic/_107_ ), .ZN(\malu/Logic/_088_ ) );
NAND2_X1 \malu/Logic/_218_ ( .A1(\malu/Logic/_057_ ), .A2(\malu/Logic/_025_ ), .ZN(\malu/Logic/_110_ ) );
AOI21_X1 \malu/Logic/_219_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_110_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_111_ ) );
AOI21_X1 \malu/Logic/_220_ ( .A(\malu/Logic/_025_ ), .B1(\malu/Logic/_100_ ), .B2(\malu/Logic/_057_ ), .ZN(\malu/Logic/_112_ ) );
OAI22_X1 \malu/Logic/_221_ ( .A1(\malu/Logic/_111_ ), .A2(\malu/Logic/_112_ ), .B1(\malu/Logic/_106_ ), .B2(\malu/Logic/_110_ ), .ZN(\malu/Logic/_091_ ) );
NAND2_X1 \malu/Logic/_222_ ( .A1(\malu/Logic/_058_ ), .A2(\malu/Logic/_026_ ), .ZN(\malu/Logic/_113_ ) );
AOI21_X1 \malu/Logic/_223_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_113_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_114_ ) );
AOI21_X1 \malu/Logic/_224_ ( .A(\malu/Logic/_026_ ), .B1(\malu/Logic/_100_ ), .B2(\malu/Logic/_058_ ), .ZN(\malu/Logic/_115_ ) );
OAI22_X1 \malu/Logic/_225_ ( .A1(\malu/Logic/_114_ ), .A2(\malu/Logic/_115_ ), .B1(\malu/Logic/_106_ ), .B2(\malu/Logic/_113_ ), .ZN(\malu/Logic/_092_ ) );
NAND2_X1 \malu/Logic/_226_ ( .A1(\malu/Logic/_059_ ), .A2(\malu/Logic/_027_ ), .ZN(\malu/Logic/_116_ ) );
AOI21_X1 \malu/Logic/_227_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_116_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_117_ ) );
AOI21_X1 \malu/Logic/_228_ ( .A(\malu/Logic/_027_ ), .B1(\malu/Logic/_100_ ), .B2(\malu/Logic/_059_ ), .ZN(\malu/Logic/_118_ ) );
OAI22_X1 \malu/Logic/_229_ ( .A1(\malu/Logic/_117_ ), .A2(\malu/Logic/_118_ ), .B1(\malu/Logic/_106_ ), .B2(\malu/Logic/_116_ ), .ZN(\malu/Logic/_093_ ) );
NAND2_X1 \malu/Logic/_230_ ( .A1(\malu/Logic/_060_ ), .A2(\malu/Logic/_028_ ), .ZN(\malu/Logic/_119_ ) );
AOI21_X1 \malu/Logic/_231_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_119_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_120_ ) );
AOI21_X1 \malu/Logic/_232_ ( .A(\malu/Logic/_028_ ), .B1(\malu/Logic/_100_ ), .B2(\malu/Logic/_060_ ), .ZN(\malu/Logic/_121_ ) );
OAI22_X1 \malu/Logic/_233_ ( .A1(\malu/Logic/_120_ ), .A2(\malu/Logic/_121_ ), .B1(\malu/Logic/_106_ ), .B2(\malu/Logic/_119_ ), .ZN(\malu/Logic/_094_ ) );
NAND2_X1 \malu/Logic/_234_ ( .A1(\malu/Logic/_061_ ), .A2(\malu/Logic/_029_ ), .ZN(\malu/Logic/_122_ ) );
AOI21_X1 \malu/Logic/_235_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_122_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_123_ ) );
AOI21_X1 \malu/Logic/_236_ ( .A(\malu/Logic/_029_ ), .B1(\malu/Logic/_100_ ), .B2(\malu/Logic/_061_ ), .ZN(\malu/Logic/_124_ ) );
OAI22_X1 \malu/Logic/_237_ ( .A1(\malu/Logic/_123_ ), .A2(\malu/Logic/_124_ ), .B1(\malu/Logic/_106_ ), .B2(\malu/Logic/_122_ ), .ZN(\malu/Logic/_095_ ) );
NAND2_X1 \malu/Logic/_238_ ( .A1(\malu/Logic/_062_ ), .A2(\malu/Logic/_030_ ), .ZN(\malu/Logic/_125_ ) );
AOI21_X1 \malu/Logic/_239_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_125_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_126_ ) );
AOI21_X1 \malu/Logic/_240_ ( .A(\malu/Logic/_030_ ), .B1(\malu/Logic/_100_ ), .B2(\malu/Logic/_062_ ), .ZN(\malu/Logic/_127_ ) );
OAI22_X1 \malu/Logic/_241_ ( .A1(\malu/Logic/_126_ ), .A2(\malu/Logic/_127_ ), .B1(\malu/Logic/_106_ ), .B2(\malu/Logic/_125_ ), .ZN(\malu/Logic/_096_ ) );
NAND2_X1 \malu/Logic/_242_ ( .A1(\malu/Logic/_063_ ), .A2(\malu/Logic/_031_ ), .ZN(\malu/Logic/_128_ ) );
AOI21_X1 \malu/Logic/_243_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_128_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_129_ ) );
AOI21_X1 \malu/Logic/_244_ ( .A(\malu/Logic/_031_ ), .B1(\malu/Logic/_100_ ), .B2(\malu/Logic/_063_ ), .ZN(\malu/Logic/_130_ ) );
OAI22_X1 \malu/Logic/_245_ ( .A1(\malu/Logic/_129_ ), .A2(\malu/Logic/_130_ ), .B1(\malu/Logic/_106_ ), .B2(\malu/Logic/_128_ ), .ZN(\malu/Logic/_097_ ) );
NAND2_X1 \malu/Logic/_246_ ( .A1(\malu/Logic/_033_ ), .A2(\malu/Logic/_001_ ), .ZN(\malu/Logic/_131_ ) );
AOI21_X1 \malu/Logic/_247_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_131_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_132_ ) );
BUF_X4 \malu/Logic/_248_ ( .A(\malu/Logic/_099_ ), .Z(\malu/Logic/_133_ ) );
AOI21_X1 \malu/Logic/_249_ ( .A(\malu/Logic/_001_ ), .B1(\malu/Logic/_133_ ), .B2(\malu/Logic/_033_ ), .ZN(\malu/Logic/_134_ ) );
OAI22_X1 \malu/Logic/_250_ ( .A1(\malu/Logic/_132_ ), .A2(\malu/Logic/_134_ ), .B1(\malu/Logic/_106_ ), .B2(\malu/Logic/_131_ ), .ZN(\malu/Logic/_067_ ) );
NAND2_X1 \malu/Logic/_251_ ( .A1(\malu/Logic/_034_ ), .A2(\malu/Logic/_002_ ), .ZN(\malu/Logic/_135_ ) );
AOI21_X1 \malu/Logic/_252_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_135_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_136_ ) );
AOI21_X1 \malu/Logic/_253_ ( .A(\malu/Logic/_002_ ), .B1(\malu/Logic/_133_ ), .B2(\malu/Logic/_034_ ), .ZN(\malu/Logic/_137_ ) );
BUF_X4 \malu/Logic/_254_ ( .A(\malu/Logic/_102_ ), .Z(\malu/Logic/_138_ ) );
OAI22_X1 \malu/Logic/_255_ ( .A1(\malu/Logic/_136_ ), .A2(\malu/Logic/_137_ ), .B1(\malu/Logic/_138_ ), .B2(\malu/Logic/_135_ ), .ZN(\malu/Logic/_068_ ) );
NAND2_X1 \malu/Logic/_256_ ( .A1(\malu/Logic/_035_ ), .A2(\malu/Logic/_003_ ), .ZN(\malu/Logic/_139_ ) );
AOI21_X1 \malu/Logic/_257_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_139_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_140_ ) );
AOI21_X1 \malu/Logic/_258_ ( .A(\malu/Logic/_003_ ), .B1(\malu/Logic/_133_ ), .B2(\malu/Logic/_035_ ), .ZN(\malu/Logic/_141_ ) );
OAI22_X1 \malu/Logic/_259_ ( .A1(\malu/Logic/_140_ ), .A2(\malu/Logic/_141_ ), .B1(\malu/Logic/_138_ ), .B2(\malu/Logic/_139_ ), .ZN(\malu/Logic/_069_ ) );
NAND2_X1 \malu/Logic/_260_ ( .A1(\malu/Logic/_036_ ), .A2(\malu/Logic/_004_ ), .ZN(\malu/Logic/_142_ ) );
AOI21_X1 \malu/Logic/_261_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_142_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_143_ ) );
AOI21_X1 \malu/Logic/_262_ ( .A(\malu/Logic/_004_ ), .B1(\malu/Logic/_133_ ), .B2(\malu/Logic/_036_ ), .ZN(\malu/Logic/_144_ ) );
OAI22_X1 \malu/Logic/_263_ ( .A1(\malu/Logic/_143_ ), .A2(\malu/Logic/_144_ ), .B1(\malu/Logic/_138_ ), .B2(\malu/Logic/_142_ ), .ZN(\malu/Logic/_070_ ) );
NAND2_X1 \malu/Logic/_264_ ( .A1(\malu/Logic/_037_ ), .A2(\malu/Logic/_005_ ), .ZN(\malu/Logic/_145_ ) );
AOI21_X1 \malu/Logic/_265_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_145_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_146_ ) );
AOI21_X1 \malu/Logic/_266_ ( .A(\malu/Logic/_005_ ), .B1(\malu/Logic/_133_ ), .B2(\malu/Logic/_037_ ), .ZN(\malu/Logic/_147_ ) );
OAI22_X1 \malu/Logic/_267_ ( .A1(\malu/Logic/_146_ ), .A2(\malu/Logic/_147_ ), .B1(\malu/Logic/_138_ ), .B2(\malu/Logic/_145_ ), .ZN(\malu/Logic/_071_ ) );
NAND2_X1 \malu/Logic/_268_ ( .A1(\malu/Logic/_038_ ), .A2(\malu/Logic/_006_ ), .ZN(\malu/Logic/_148_ ) );
AOI21_X1 \malu/Logic/_269_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_148_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_149_ ) );
AOI21_X1 \malu/Logic/_270_ ( .A(\malu/Logic/_006_ ), .B1(\malu/Logic/_133_ ), .B2(\malu/Logic/_038_ ), .ZN(\malu/Logic/_150_ ) );
OAI22_X1 \malu/Logic/_271_ ( .A1(\malu/Logic/_149_ ), .A2(\malu/Logic/_150_ ), .B1(\malu/Logic/_138_ ), .B2(\malu/Logic/_148_ ), .ZN(\malu/Logic/_072_ ) );
NAND2_X1 \malu/Logic/_272_ ( .A1(\malu/Logic/_039_ ), .A2(\malu/Logic/_007_ ), .ZN(\malu/Logic/_151_ ) );
AOI21_X1 \malu/Logic/_273_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_151_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_152_ ) );
AOI21_X1 \malu/Logic/_274_ ( .A(\malu/Logic/_007_ ), .B1(\malu/Logic/_133_ ), .B2(\malu/Logic/_039_ ), .ZN(\malu/Logic/_153_ ) );
OAI22_X1 \malu/Logic/_275_ ( .A1(\malu/Logic/_152_ ), .A2(\malu/Logic/_153_ ), .B1(\malu/Logic/_138_ ), .B2(\malu/Logic/_151_ ), .ZN(\malu/Logic/_073_ ) );
NAND2_X1 \malu/Logic/_276_ ( .A1(\malu/Logic/_040_ ), .A2(\malu/Logic/_008_ ), .ZN(\malu/Logic/_154_ ) );
AOI21_X1 \malu/Logic/_277_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_154_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_155_ ) );
AOI21_X1 \malu/Logic/_278_ ( .A(\malu/Logic/_008_ ), .B1(\malu/Logic/_133_ ), .B2(\malu/Logic/_040_ ), .ZN(\malu/Logic/_156_ ) );
OAI22_X1 \malu/Logic/_279_ ( .A1(\malu/Logic/_155_ ), .A2(\malu/Logic/_156_ ), .B1(\malu/Logic/_138_ ), .B2(\malu/Logic/_154_ ), .ZN(\malu/Logic/_074_ ) );
NAND2_X1 \malu/Logic/_280_ ( .A1(\malu/Logic/_041_ ), .A2(\malu/Logic/_009_ ), .ZN(\malu/Logic/_157_ ) );
AOI21_X1 \malu/Logic/_281_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_157_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_158_ ) );
AOI21_X1 \malu/Logic/_282_ ( .A(\malu/Logic/_009_ ), .B1(\malu/Logic/_133_ ), .B2(\malu/Logic/_041_ ), .ZN(\malu/Logic/_159_ ) );
OAI22_X1 \malu/Logic/_283_ ( .A1(\malu/Logic/_158_ ), .A2(\malu/Logic/_159_ ), .B1(\malu/Logic/_138_ ), .B2(\malu/Logic/_157_ ), .ZN(\malu/Logic/_075_ ) );
NAND2_X1 \malu/Logic/_284_ ( .A1(\malu/Logic/_042_ ), .A2(\malu/Logic/_010_ ), .ZN(\malu/Logic/_160_ ) );
AOI21_X1 \malu/Logic/_285_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_160_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_161_ ) );
AOI21_X1 \malu/Logic/_286_ ( .A(\malu/Logic/_010_ ), .B1(\malu/Logic/_133_ ), .B2(\malu/Logic/_042_ ), .ZN(\malu/Logic/_162_ ) );
OAI22_X1 \malu/Logic/_287_ ( .A1(\malu/Logic/_161_ ), .A2(\malu/Logic/_162_ ), .B1(\malu/Logic/_138_ ), .B2(\malu/Logic/_160_ ), .ZN(\malu/Logic/_076_ ) );
NAND2_X1 \malu/Logic/_288_ ( .A1(\malu/Logic/_044_ ), .A2(\malu/Logic/_012_ ), .ZN(\malu/Logic/_163_ ) );
AOI21_X1 \malu/Logic/_289_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_163_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_164_ ) );
BUF_X4 \malu/Logic/_290_ ( .A(\malu/Logic/_099_ ), .Z(\malu/Logic/_165_ ) );
AOI21_X1 \malu/Logic/_291_ ( .A(\malu/Logic/_012_ ), .B1(\malu/Logic/_165_ ), .B2(\malu/Logic/_044_ ), .ZN(\malu/Logic/_166_ ) );
OAI22_X1 \malu/Logic/_292_ ( .A1(\malu/Logic/_164_ ), .A2(\malu/Logic/_166_ ), .B1(\malu/Logic/_138_ ), .B2(\malu/Logic/_163_ ), .ZN(\malu/Logic/_078_ ) );
NAND2_X1 \malu/Logic/_293_ ( .A1(\malu/Logic/_045_ ), .A2(\malu/Logic/_013_ ), .ZN(\malu/Logic/_167_ ) );
AOI21_X1 \malu/Logic/_294_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_167_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_168_ ) );
AOI21_X1 \malu/Logic/_295_ ( .A(\malu/Logic/_013_ ), .B1(\malu/Logic/_165_ ), .B2(\malu/Logic/_045_ ), .ZN(\malu/Logic/_169_ ) );
BUF_X4 \malu/Logic/_296_ ( .A(\malu/Logic/_102_ ), .Z(\malu/Logic/_170_ ) );
OAI22_X1 \malu/Logic/_297_ ( .A1(\malu/Logic/_168_ ), .A2(\malu/Logic/_169_ ), .B1(\malu/Logic/_170_ ), .B2(\malu/Logic/_167_ ), .ZN(\malu/Logic/_079_ ) );
NAND2_X1 \malu/Logic/_298_ ( .A1(\malu/Logic/_046_ ), .A2(\malu/Logic/_014_ ), .ZN(\malu/Logic/_171_ ) );
AOI21_X1 \malu/Logic/_299_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_171_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_172_ ) );
AOI21_X1 \malu/Logic/_300_ ( .A(\malu/Logic/_014_ ), .B1(\malu/Logic/_165_ ), .B2(\malu/Logic/_046_ ), .ZN(\malu/Logic/_173_ ) );
OAI22_X1 \malu/Logic/_301_ ( .A1(\malu/Logic/_172_ ), .A2(\malu/Logic/_173_ ), .B1(\malu/Logic/_170_ ), .B2(\malu/Logic/_171_ ), .ZN(\malu/Logic/_080_ ) );
NAND2_X1 \malu/Logic/_302_ ( .A1(\malu/Logic/_047_ ), .A2(\malu/Logic/_015_ ), .ZN(\malu/Logic/_174_ ) );
AOI21_X1 \malu/Logic/_303_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_174_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_175_ ) );
AOI21_X1 \malu/Logic/_304_ ( .A(\malu/Logic/_015_ ), .B1(\malu/Logic/_165_ ), .B2(\malu/Logic/_047_ ), .ZN(\malu/Logic/_176_ ) );
OAI22_X1 \malu/Logic/_305_ ( .A1(\malu/Logic/_175_ ), .A2(\malu/Logic/_176_ ), .B1(\malu/Logic/_170_ ), .B2(\malu/Logic/_174_ ), .ZN(\malu/Logic/_081_ ) );
NAND2_X1 \malu/Logic/_306_ ( .A1(\malu/Logic/_048_ ), .A2(\malu/Logic/_016_ ), .ZN(\malu/Logic/_177_ ) );
AOI21_X1 \malu/Logic/_307_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_177_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_178_ ) );
AOI21_X1 \malu/Logic/_308_ ( .A(\malu/Logic/_016_ ), .B1(\malu/Logic/_165_ ), .B2(\malu/Logic/_048_ ), .ZN(\malu/Logic/_179_ ) );
OAI22_X1 \malu/Logic/_309_ ( .A1(\malu/Logic/_178_ ), .A2(\malu/Logic/_179_ ), .B1(\malu/Logic/_170_ ), .B2(\malu/Logic/_177_ ), .ZN(\malu/Logic/_082_ ) );
NAND2_X1 \malu/Logic/_310_ ( .A1(\malu/Logic/_049_ ), .A2(\malu/Logic/_017_ ), .ZN(\malu/Logic/_180_ ) );
AOI21_X1 \malu/Logic/_311_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_180_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_181_ ) );
AOI21_X2 \malu/Logic/_312_ ( .A(\malu/Logic/_017_ ), .B1(\malu/Logic/_165_ ), .B2(\malu/Logic/_049_ ), .ZN(\malu/Logic/_182_ ) );
OAI22_X1 \malu/Logic/_313_ ( .A1(\malu/Logic/_181_ ), .A2(\malu/Logic/_182_ ), .B1(\malu/Logic/_170_ ), .B2(\malu/Logic/_180_ ), .ZN(\malu/Logic/_083_ ) );
NAND2_X1 \malu/Logic/_314_ ( .A1(\malu/Logic/_050_ ), .A2(\malu/Logic/_018_ ), .ZN(\malu/Logic/_183_ ) );
AOI21_X1 \malu/Logic/_315_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_183_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_184_ ) );
AOI21_X2 \malu/Logic/_316_ ( .A(\malu/Logic/_018_ ), .B1(\malu/Logic/_165_ ), .B2(\malu/Logic/_050_ ), .ZN(\malu/Logic/_185_ ) );
OAI22_X1 \malu/Logic/_317_ ( .A1(\malu/Logic/_184_ ), .A2(\malu/Logic/_185_ ), .B1(\malu/Logic/_170_ ), .B2(\malu/Logic/_183_ ), .ZN(\malu/Logic/_084_ ) );
NAND2_X1 \malu/Logic/_318_ ( .A1(\malu/Logic/_051_ ), .A2(\malu/Logic/_019_ ), .ZN(\malu/Logic/_186_ ) );
AOI21_X1 \malu/Logic/_319_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_186_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_187_ ) );
AOI21_X2 \malu/Logic/_320_ ( .A(\malu/Logic/_019_ ), .B1(\malu/Logic/_165_ ), .B2(\malu/Logic/_051_ ), .ZN(\malu/Logic/_188_ ) );
OAI22_X1 \malu/Logic/_321_ ( .A1(\malu/Logic/_187_ ), .A2(\malu/Logic/_188_ ), .B1(\malu/Logic/_170_ ), .B2(\malu/Logic/_186_ ), .ZN(\malu/Logic/_085_ ) );
NAND2_X1 \malu/Logic/_322_ ( .A1(\malu/Logic/_052_ ), .A2(\malu/Logic/_020_ ), .ZN(\malu/Logic/_189_ ) );
AOI21_X1 \malu/Logic/_323_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_189_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_190_ ) );
AOI21_X2 \malu/Logic/_324_ ( .A(\malu/Logic/_020_ ), .B1(\malu/Logic/_165_ ), .B2(\malu/Logic/_052_ ), .ZN(\malu/Logic/_191_ ) );
OAI22_X1 \malu/Logic/_325_ ( .A1(\malu/Logic/_190_ ), .A2(\malu/Logic/_191_ ), .B1(\malu/Logic/_170_ ), .B2(\malu/Logic/_189_ ), .ZN(\malu/Logic/_086_ ) );
NAND2_X1 \malu/Logic/_326_ ( .A1(\malu/Logic/_053_ ), .A2(\malu/Logic/_021_ ), .ZN(\malu/Logic/_192_ ) );
AOI21_X1 \malu/Logic/_327_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_192_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_193_ ) );
AOI21_X1 \malu/Logic/_328_ ( .A(\malu/Logic/_021_ ), .B1(\malu/Logic/_165_ ), .B2(\malu/Logic/_053_ ), .ZN(\malu/Logic/_194_ ) );
OAI22_X1 \malu/Logic/_329_ ( .A1(\malu/Logic/_193_ ), .A2(\malu/Logic/_194_ ), .B1(\malu/Logic/_170_ ), .B2(\malu/Logic/_192_ ), .ZN(\malu/Logic/_087_ ) );
NAND2_X1 \malu/Logic/_330_ ( .A1(\malu/Logic/_055_ ), .A2(\malu/Logic/_023_ ), .ZN(\malu/Logic/_195_ ) );
AOI21_X1 \malu/Logic/_331_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_195_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_196_ ) );
AOI21_X1 \malu/Logic/_332_ ( .A(\malu/Logic/_023_ ), .B1(\malu/Logic/_099_ ), .B2(\malu/Logic/_055_ ), .ZN(\malu/Logic/_197_ ) );
OAI22_X1 \malu/Logic/_333_ ( .A1(\malu/Logic/_196_ ), .A2(\malu/Logic/_197_ ), .B1(\malu/Logic/_170_ ), .B2(\malu/Logic/_195_ ), .ZN(\malu/Logic/_089_ ) );
NAND2_X1 \malu/Logic/_334_ ( .A1(\malu/Logic/_056_ ), .A2(\malu/Logic/_024_ ), .ZN(\malu/Logic/_198_ ) );
AOI21_X1 \malu/Logic/_335_ ( .A(\malu/Logic/_064_ ), .B1(\malu/Logic/_198_ ), .B2(\malu/Logic/_065_ ), .ZN(\malu/Logic/_199_ ) );
AOI21_X1 \malu/Logic/_336_ ( .A(\malu/Logic/_024_ ), .B1(\malu/Logic/_099_ ), .B2(\malu/Logic/_056_ ), .ZN(\malu/Logic/_200_ ) );
OAI22_X1 \malu/Logic/_337_ ( .A1(\malu/Logic/_199_ ), .A2(\malu/Logic/_200_ ), .B1(\malu/Logic/_102_ ), .B2(\malu/Logic/_198_ ), .ZN(\malu/Logic/_090_ ) );
BUF_X1 \malu/Logic/_338_ ( .A(\alu_b[0] ), .Z(\malu/Logic/_032_ ) );
BUF_X1 \malu/Logic/_339_ ( .A(\alu_a[0] ), .Z(\malu/Logic/_000_ ) );
BUF_X1 \malu/Logic/_340_ ( .A(\malu/logic_ctl[0] ), .Z(\malu/Logic/_064_ ) );
BUF_X1 \malu/Logic/_341_ ( .A(\malu/logic_ctl[1] ), .Z(\malu/Logic/_065_ ) );
BUF_X1 \malu/Logic/_342_ ( .A(\malu/Logic/_066_ ), .Z(\malu/logic_result[0] ) );
BUF_X1 \malu/Logic/_343_ ( .A(\alu_b[1] ), .Z(\malu/Logic/_043_ ) );
BUF_X1 \malu/Logic/_344_ ( .A(\alu_a[1] ), .Z(\malu/Logic/_011_ ) );
BUF_X1 \malu/Logic/_345_ ( .A(\malu/Logic/_077_ ), .Z(\malu/logic_result[1] ) );
BUF_X1 \malu/Logic/_346_ ( .A(\alu_b[2] ), .Z(\malu/Logic/_054_ ) );
BUF_X1 \malu/Logic/_347_ ( .A(\alu_a[2] ), .Z(\malu/Logic/_022_ ) );
BUF_X1 \malu/Logic/_348_ ( .A(\malu/Logic/_088_ ), .Z(\malu/logic_result[2] ) );
BUF_X1 \malu/Logic/_349_ ( .A(\alu_b[3] ), .Z(\malu/Logic/_057_ ) );
BUF_X1 \malu/Logic/_350_ ( .A(\alu_a[3] ), .Z(\malu/Logic/_025_ ) );
BUF_X1 \malu/Logic/_351_ ( .A(\malu/Logic/_091_ ), .Z(\malu/logic_result[3] ) );
BUF_X1 \malu/Logic/_352_ ( .A(\alu_b[4] ), .Z(\malu/Logic/_058_ ) );
BUF_X1 \malu/Logic/_353_ ( .A(\alu_a[4] ), .Z(\malu/Logic/_026_ ) );
BUF_X1 \malu/Logic/_354_ ( .A(\malu/Logic/_092_ ), .Z(\malu/logic_result[4] ) );
BUF_X1 \malu/Logic/_355_ ( .A(\alu_b[5] ), .Z(\malu/Logic/_059_ ) );
BUF_X1 \malu/Logic/_356_ ( .A(\alu_a[5] ), .Z(\malu/Logic/_027_ ) );
BUF_X1 \malu/Logic/_357_ ( .A(\malu/Logic/_093_ ), .Z(\malu/logic_result[5] ) );
BUF_X1 \malu/Logic/_358_ ( .A(\alu_b[6] ), .Z(\malu/Logic/_060_ ) );
BUF_X1 \malu/Logic/_359_ ( .A(\alu_a[6] ), .Z(\malu/Logic/_028_ ) );
BUF_X1 \malu/Logic/_360_ ( .A(\malu/Logic/_094_ ), .Z(\malu/logic_result[6] ) );
BUF_X1 \malu/Logic/_361_ ( .A(\alu_b[7] ), .Z(\malu/Logic/_061_ ) );
BUF_X1 \malu/Logic/_362_ ( .A(\alu_a[7] ), .Z(\malu/Logic/_029_ ) );
BUF_X1 \malu/Logic/_363_ ( .A(\malu/Logic/_095_ ), .Z(\malu/logic_result[7] ) );
BUF_X1 \malu/Logic/_364_ ( .A(\alu_b[8] ), .Z(\malu/Logic/_062_ ) );
BUF_X1 \malu/Logic/_365_ ( .A(\alu_a[8] ), .Z(\malu/Logic/_030_ ) );
BUF_X1 \malu/Logic/_366_ ( .A(\malu/Logic/_096_ ), .Z(\malu/logic_result[8] ) );
BUF_X1 \malu/Logic/_367_ ( .A(\alu_b[9] ), .Z(\malu/Logic/_063_ ) );
BUF_X1 \malu/Logic/_368_ ( .A(\alu_a[9] ), .Z(\malu/Logic/_031_ ) );
BUF_X1 \malu/Logic/_369_ ( .A(\malu/Logic/_097_ ), .Z(\malu/logic_result[9] ) );
BUF_X1 \malu/Logic/_370_ ( .A(\alu_b[10] ), .Z(\malu/Logic/_033_ ) );
BUF_X1 \malu/Logic/_371_ ( .A(\alu_a[10] ), .Z(\malu/Logic/_001_ ) );
BUF_X1 \malu/Logic/_372_ ( .A(\malu/Logic/_067_ ), .Z(\malu/logic_result[10] ) );
BUF_X1 \malu/Logic/_373_ ( .A(\alu_b[11] ), .Z(\malu/Logic/_034_ ) );
BUF_X1 \malu/Logic/_374_ ( .A(\alu_a[11] ), .Z(\malu/Logic/_002_ ) );
BUF_X1 \malu/Logic/_375_ ( .A(\malu/Logic/_068_ ), .Z(\malu/logic_result[11] ) );
BUF_X1 \malu/Logic/_376_ ( .A(\alu_b[12] ), .Z(\malu/Logic/_035_ ) );
BUF_X1 \malu/Logic/_377_ ( .A(\alu_a[12] ), .Z(\malu/Logic/_003_ ) );
BUF_X1 \malu/Logic/_378_ ( .A(\malu/Logic/_069_ ), .Z(\malu/logic_result[12] ) );
BUF_X1 \malu/Logic/_379_ ( .A(\alu_b[13] ), .Z(\malu/Logic/_036_ ) );
BUF_X1 \malu/Logic/_380_ ( .A(\alu_a[13] ), .Z(\malu/Logic/_004_ ) );
BUF_X1 \malu/Logic/_381_ ( .A(\malu/Logic/_070_ ), .Z(\malu/logic_result[13] ) );
BUF_X1 \malu/Logic/_382_ ( .A(\alu_b[14] ), .Z(\malu/Logic/_037_ ) );
BUF_X1 \malu/Logic/_383_ ( .A(\alu_a[14] ), .Z(\malu/Logic/_005_ ) );
BUF_X1 \malu/Logic/_384_ ( .A(\malu/Logic/_071_ ), .Z(\malu/logic_result[14] ) );
BUF_X1 \malu/Logic/_385_ ( .A(\alu_b[15] ), .Z(\malu/Logic/_038_ ) );
BUF_X1 \malu/Logic/_386_ ( .A(\alu_a[15] ), .Z(\malu/Logic/_006_ ) );
BUF_X1 \malu/Logic/_387_ ( .A(\malu/Logic/_072_ ), .Z(\malu/logic_result[15] ) );
BUF_X1 \malu/Logic/_388_ ( .A(\alu_b[16] ), .Z(\malu/Logic/_039_ ) );
BUF_X1 \malu/Logic/_389_ ( .A(\alu_a[16] ), .Z(\malu/Logic/_007_ ) );
BUF_X1 \malu/Logic/_390_ ( .A(\malu/Logic/_073_ ), .Z(\malu/logic_result[16] ) );
BUF_X1 \malu/Logic/_391_ ( .A(\alu_b[17] ), .Z(\malu/Logic/_040_ ) );
BUF_X1 \malu/Logic/_392_ ( .A(\alu_a[17] ), .Z(\malu/Logic/_008_ ) );
BUF_X1 \malu/Logic/_393_ ( .A(\malu/Logic/_074_ ), .Z(\malu/logic_result[17] ) );
BUF_X1 \malu/Logic/_394_ ( .A(\alu_b[18] ), .Z(\malu/Logic/_041_ ) );
BUF_X1 \malu/Logic/_395_ ( .A(\alu_a[18] ), .Z(\malu/Logic/_009_ ) );
BUF_X1 \malu/Logic/_396_ ( .A(\malu/Logic/_075_ ), .Z(\malu/logic_result[18] ) );
BUF_X1 \malu/Logic/_397_ ( .A(\alu_b[19] ), .Z(\malu/Logic/_042_ ) );
BUF_X1 \malu/Logic/_398_ ( .A(\alu_a[19] ), .Z(\malu/Logic/_010_ ) );
BUF_X1 \malu/Logic/_399_ ( .A(\malu/Logic/_076_ ), .Z(\malu/logic_result[19] ) );
BUF_X1 \malu/Logic/_400_ ( .A(\alu_b[20] ), .Z(\malu/Logic/_044_ ) );
BUF_X1 \malu/Logic/_401_ ( .A(\alu_a[20] ), .Z(\malu/Logic/_012_ ) );
BUF_X1 \malu/Logic/_402_ ( .A(\malu/Logic/_078_ ), .Z(\malu/logic_result[20] ) );
BUF_X1 \malu/Logic/_403_ ( .A(\alu_b[21] ), .Z(\malu/Logic/_045_ ) );
BUF_X1 \malu/Logic/_404_ ( .A(\alu_a[21] ), .Z(\malu/Logic/_013_ ) );
BUF_X1 \malu/Logic/_405_ ( .A(\malu/Logic/_079_ ), .Z(\malu/logic_result[21] ) );
BUF_X1 \malu/Logic/_406_ ( .A(\alu_b[22] ), .Z(\malu/Logic/_046_ ) );
BUF_X1 \malu/Logic/_407_ ( .A(\alu_a[22] ), .Z(\malu/Logic/_014_ ) );
BUF_X1 \malu/Logic/_408_ ( .A(\malu/Logic/_080_ ), .Z(\malu/logic_result[22] ) );
BUF_X1 \malu/Logic/_409_ ( .A(\alu_b[23] ), .Z(\malu/Logic/_047_ ) );
BUF_X1 \malu/Logic/_410_ ( .A(\alu_a[23] ), .Z(\malu/Logic/_015_ ) );
BUF_X1 \malu/Logic/_411_ ( .A(\malu/Logic/_081_ ), .Z(\malu/logic_result[23] ) );
BUF_X1 \malu/Logic/_412_ ( .A(\alu_b[24] ), .Z(\malu/Logic/_048_ ) );
BUF_X1 \malu/Logic/_413_ ( .A(\alu_a[24] ), .Z(\malu/Logic/_016_ ) );
BUF_X1 \malu/Logic/_414_ ( .A(\malu/Logic/_082_ ), .Z(\malu/logic_result[24] ) );
BUF_X1 \malu/Logic/_415_ ( .A(\alu_b[25] ), .Z(\malu/Logic/_049_ ) );
BUF_X1 \malu/Logic/_416_ ( .A(\alu_a[25] ), .Z(\malu/Logic/_017_ ) );
BUF_X1 \malu/Logic/_417_ ( .A(\malu/Logic/_083_ ), .Z(\malu/logic_result[25] ) );
BUF_X1 \malu/Logic/_418_ ( .A(\alu_b[26] ), .Z(\malu/Logic/_050_ ) );
BUF_X1 \malu/Logic/_419_ ( .A(\alu_a[26] ), .Z(\malu/Logic/_018_ ) );
BUF_X1 \malu/Logic/_420_ ( .A(\malu/Logic/_084_ ), .Z(\malu/logic_result[26] ) );
BUF_X1 \malu/Logic/_421_ ( .A(\alu_b[27] ), .Z(\malu/Logic/_051_ ) );
BUF_X1 \malu/Logic/_422_ ( .A(\alu_a[27] ), .Z(\malu/Logic/_019_ ) );
BUF_X1 \malu/Logic/_423_ ( .A(\malu/Logic/_085_ ), .Z(\malu/logic_result[27] ) );
BUF_X1 \malu/Logic/_424_ ( .A(\alu_b[28] ), .Z(\malu/Logic/_052_ ) );
BUF_X1 \malu/Logic/_425_ ( .A(\alu_a[28] ), .Z(\malu/Logic/_020_ ) );
BUF_X1 \malu/Logic/_426_ ( .A(\malu/Logic/_086_ ), .Z(\malu/logic_result[28] ) );
BUF_X1 \malu/Logic/_427_ ( .A(\alu_b[29] ), .Z(\malu/Logic/_053_ ) );
BUF_X1 \malu/Logic/_428_ ( .A(\alu_a[29] ), .Z(\malu/Logic/_021_ ) );
BUF_X1 \malu/Logic/_429_ ( .A(\malu/Logic/_087_ ), .Z(\malu/logic_result[29] ) );
BUF_X1 \malu/Logic/_430_ ( .A(\alu_b[30] ), .Z(\malu/Logic/_055_ ) );
BUF_X1 \malu/Logic/_431_ ( .A(\alu_a[30] ), .Z(\malu/Logic/_023_ ) );
BUF_X1 \malu/Logic/_432_ ( .A(\malu/Logic/_089_ ), .Z(\malu/logic_result[30] ) );
BUF_X1 \malu/Logic/_433_ ( .A(\alu_b[31] ), .Z(\malu/Logic/_056_ ) );
BUF_X1 \malu/Logic/_434_ ( .A(\alu_a[31] ), .Z(\malu/Logic/_024_ ) );
BUF_X1 \malu/Logic/_435_ ( .A(\malu/Logic/_090_ ), .Z(\malu/logic_result[31] ) );
AND2_X2 \malu/Shift/_0753_ ( .A1(\malu/Shift/_0714_ ), .A2(\malu/Shift/_0715_ ), .ZN(\malu/Shift/_0635_ ) );
NOR2_X1 \malu/Shift/_0754_ ( .A1(\malu/Shift/_0714_ ), .A2(\malu/Shift/_0715_ ), .ZN(\malu/Shift/_0646_ ) );
NOR2_X1 \malu/Shift/_0755_ ( .A1(\malu/Shift/_0635_ ), .A2(\malu/Shift/_0646_ ), .ZN(\malu/Shift/_0656_ ) );
INV_X1 \malu/Shift/_0756_ ( .A(\malu/Shift/_0001_ ), .ZN(\malu/Shift/_0666_ ) );
NOR2_X1 \malu/Shift/_0757_ ( .A1(\malu/Shift/_0666_ ), .A2(\malu/Shift/_0716_ ), .ZN(\malu/Shift/_0676_ ) );
AND2_X4 \malu/Shift/_0758_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0002_ ), .ZN(\malu/Shift/_0686_ ) );
INV_X32 \malu/Shift/_0759_ ( .A(\malu/Shift/_0717_ ), .ZN(\malu/Shift/_0692_ ) );
BUF_X8 \malu/Shift/_0760_ ( .A(\malu/Shift/_0692_ ), .Z(\malu/Shift/_0693_ ) );
OR3_X4 \malu/Shift/_0761_ ( .A1(\malu/Shift/_0676_ ), .A2(\malu/Shift/_0686_ ), .A3(\malu/Shift/_0693_ ), .ZN(\malu/Shift/_0694_ ) );
INV_X1 \malu/Shift/_0762_ ( .A(\malu/Shift/_0030_ ), .ZN(\malu/Shift/_0695_ ) );
NOR2_X1 \malu/Shift/_0763_ ( .A1(\malu/Shift/_0695_ ), .A2(\malu/Shift/_0716_ ), .ZN(\malu/Shift/_0696_ ) );
AND2_X4 \malu/Shift/_0764_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0031_ ), .ZN(\malu/Shift/_0697_ ) );
OR3_X2 \malu/Shift/_0765_ ( .A1(\malu/Shift/_0696_ ), .A2(\malu/Shift/_0697_ ), .A3(\malu/Shift/_0717_ ), .ZN(\malu/Shift/_0698_ ) );
AOI21_X1 \malu/Shift/_0766_ ( .A(\malu/Shift/_0718_ ), .B1(\malu/Shift/_0694_ ), .B2(\malu/Shift/_0698_ ), .ZN(\malu/Shift/_0699_ ) );
BUF_X4 \malu/Shift/_0767_ ( .A(\malu/Shift/_0692_ ), .Z(\malu/Shift/_0700_ ) );
INV_X1 \malu/Shift/_0768_ ( .A(\malu/Shift/_0003_ ), .ZN(\malu/Shift/_0701_ ) );
NOR2_X1 \malu/Shift/_0769_ ( .A1(\malu/Shift/_0701_ ), .A2(\malu/Shift/_0716_ ), .ZN(\malu/Shift/_0702_ ) );
AND2_X1 \malu/Shift/_0770_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0004_ ), .ZN(\malu/Shift/_0703_ ) );
OAI21_X1 \malu/Shift/_0771_ ( .A(\malu/Shift/_0700_ ), .B1(\malu/Shift/_0702_ ), .B2(\malu/Shift/_0703_ ), .ZN(\malu/Shift/_0704_ ) );
INV_X1 \malu/Shift/_0772_ ( .A(\malu/Shift/_0005_ ), .ZN(\malu/Shift/_0705_ ) );
NOR2_X1 \malu/Shift/_0773_ ( .A1(\malu/Shift/_0705_ ), .A2(\malu/Shift/_0716_ ), .ZN(\malu/Shift/_0706_ ) );
AND2_X1 \malu/Shift/_0774_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0006_ ), .ZN(\malu/Shift/_0707_ ) );
OAI21_X1 \malu/Shift/_0775_ ( .A(\malu/Shift/_0717_ ), .B1(\malu/Shift/_0706_ ), .B2(\malu/Shift/_0707_ ), .ZN(\malu/Shift/_0708_ ) );
AND3_X1 \malu/Shift/_0776_ ( .A1(\malu/Shift/_0704_ ), .A2(\malu/Shift/_0708_ ), .A3(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0709_ ) );
INV_X2 \malu/Shift/_0777_ ( .A(\malu/Shift/_0719_ ), .ZN(\malu/Shift/_0710_ ) );
BUF_X4 \malu/Shift/_0778_ ( .A(\malu/Shift/_0710_ ), .Z(\malu/Shift/_0711_ ) );
OR3_X1 \malu/Shift/_0779_ ( .A1(\malu/Shift/_0699_ ), .A2(\malu/Shift/_0709_ ), .A3(\malu/Shift/_0711_ ), .ZN(\malu/Shift/_0712_ ) );
INV_X1 \malu/Shift/_0780_ ( .A(\malu/Shift/_0000_ ), .ZN(\malu/Shift/_0713_ ) );
NOR2_X1 \malu/Shift/_0781_ ( .A1(\malu/Shift/_0713_ ), .A2(\malu/Shift/_0716_ ), .ZN(\malu/Shift/_0032_ ) );
BUF_X4 \malu/Shift/_0782_ ( .A(\malu/Shift/_0693_ ), .Z(\malu/Shift/_0033_ ) );
BUF_X4 \malu/Shift/_0783_ ( .A(\malu/Shift/_0033_ ), .Z(\malu/Shift/_0034_ ) );
AND2_X1 \malu/Shift/_0784_ ( .A1(\malu/Shift/_0032_ ), .A2(\malu/Shift/_0034_ ), .ZN(\malu/Shift/_0035_ ) );
INV_X1 \malu/Shift/_0785_ ( .A(\malu/Shift/_0035_ ), .ZN(\malu/Shift/_0036_ ) );
AND2_X1 \malu/Shift/_0786_ ( .A1(\malu/Shift/_0011_ ), .A2(\malu/Shift/_0716_ ), .ZN(\malu/Shift/_0037_ ) );
BUF_X2 \malu/Shift/_0787_ ( .A(\malu/Shift/_0700_ ), .Z(\malu/Shift/_0038_ ) );
BUF_X4 \malu/Shift/_0788_ ( .A(\malu/Shift/_0038_ ), .Z(\malu/Shift/_0039_ ) );
AOI21_X1 \malu/Shift/_0789_ ( .A(\malu/Shift/_0718_ ), .B1(\malu/Shift/_0037_ ), .B2(\malu/Shift/_0039_ ), .ZN(\malu/Shift/_0040_ ) );
INV_X32 \malu/Shift/_0790_ ( .A(\malu/Shift/_0716_ ), .ZN(\malu/Shift/_0041_ ) );
BUF_X32 \malu/Shift/_0791_ ( .A(\malu/Shift/_0041_ ), .Z(\malu/Shift/_0042_ ) );
AND2_X4 \malu/Shift/_0792_ ( .A1(\malu/Shift/_0042_ ), .A2(\malu/Shift/_0022_ ), .ZN(\malu/Shift/_0043_ ) );
AND2_X1 \malu/Shift/_0793_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0025_ ), .ZN(\malu/Shift/_0044_ ) );
NOR2_X1 \malu/Shift/_0794_ ( .A1(\malu/Shift/_0043_ ), .A2(\malu/Shift/_0044_ ), .ZN(\malu/Shift/_0045_ ) );
OAI211_X2 \malu/Shift/_0795_ ( .A(\malu/Shift/_0036_ ), .B(\malu/Shift/_0040_ ), .C1(\malu/Shift/_0039_ ), .C2(\malu/Shift/_0045_ ), .ZN(\malu/Shift/_0046_ ) );
BUF_X4 \malu/Shift/_0796_ ( .A(\malu/Shift/_0710_ ), .Z(\malu/Shift/_0047_ ) );
BUF_X4 \malu/Shift/_0797_ ( .A(\malu/Shift/_0047_ ), .Z(\malu/Shift/_0048_ ) );
INV_X1 \malu/Shift/_0798_ ( .A(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0049_ ) );
BUF_X4 \malu/Shift/_0799_ ( .A(\malu/Shift/_0049_ ), .Z(\malu/Shift/_0050_ ) );
BUF_X4 \malu/Shift/_0800_ ( .A(\malu/Shift/_0050_ ), .Z(\malu/Shift/_0051_ ) );
BUF_X4 \malu/Shift/_0801_ ( .A(\malu/Shift/_0051_ ), .Z(\malu/Shift/_0052_ ) );
BUF_X4 \malu/Shift/_0802_ ( .A(\malu/Shift/_0052_ ), .Z(\malu/Shift/_0053_ ) );
AND2_X4 \malu/Shift/_0803_ ( .A1(\malu/Shift/_0042_ ), .A2(\malu/Shift/_0026_ ), .ZN(\malu/Shift/_0054_ ) );
AND2_X4 \malu/Shift/_0804_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0027_ ), .ZN(\malu/Shift/_0055_ ) );
OAI21_X1 \malu/Shift/_0805_ ( .A(\malu/Shift/_0033_ ), .B1(\malu/Shift/_0054_ ), .B2(\malu/Shift/_0055_ ), .ZN(\malu/Shift/_0056_ ) );
INV_X1 \malu/Shift/_0806_ ( .A(\malu/Shift/_0028_ ), .ZN(\malu/Shift/_0057_ ) );
NOR2_X1 \malu/Shift/_0807_ ( .A1(\malu/Shift/_0057_ ), .A2(\malu/Shift/_0716_ ), .ZN(\malu/Shift/_0058_ ) );
AND2_X4 \malu/Shift/_0808_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0029_ ), .ZN(\malu/Shift/_0059_ ) );
OAI21_X1 \malu/Shift/_0809_ ( .A(\malu/Shift/_0717_ ), .B1(\malu/Shift/_0058_ ), .B2(\malu/Shift/_0059_ ), .ZN(\malu/Shift/_0060_ ) );
NAND2_X1 \malu/Shift/_0810_ ( .A1(\malu/Shift/_0056_ ), .A2(\malu/Shift/_0060_ ), .ZN(\malu/Shift/_0061_ ) );
OAI211_X2 \malu/Shift/_0811_ ( .A(\malu/Shift/_0046_ ), .B(\malu/Shift/_0048_ ), .C1(\malu/Shift/_0053_ ), .C2(\malu/Shift/_0061_ ), .ZN(\malu/Shift/_0062_ ) );
AOI21_X1 \malu/Shift/_0812_ ( .A(\malu/Shift/_0720_ ), .B1(\malu/Shift/_0712_ ), .B2(\malu/Shift/_0062_ ), .ZN(\malu/Shift/_0063_ ) );
BUF_X4 \malu/Shift/_0813_ ( .A(\malu/Shift/_0710_ ), .Z(\malu/Shift/_0064_ ) );
AND2_X1 \malu/Shift/_0814_ ( .A1(\malu/Shift/_0041_ ), .A2(\malu/Shift/_0014_ ), .ZN(\malu/Shift/_0065_ ) );
AND2_X4 \malu/Shift/_0815_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0015_ ), .ZN(\malu/Shift/_0066_ ) );
OR3_X1 \malu/Shift/_0816_ ( .A1(\malu/Shift/_0065_ ), .A2(\malu/Shift/_0066_ ), .A3(\malu/Shift/_0700_ ), .ZN(\malu/Shift/_0067_ ) );
INV_X1 \malu/Shift/_0817_ ( .A(\malu/Shift/_0012_ ), .ZN(\malu/Shift/_0068_ ) );
NOR2_X1 \malu/Shift/_0818_ ( .A1(\malu/Shift/_0068_ ), .A2(\malu/Shift/_0716_ ), .ZN(\malu/Shift/_0069_ ) );
AND2_X1 \malu/Shift/_0819_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0013_ ), .ZN(\malu/Shift/_0070_ ) );
OR3_X1 \malu/Shift/_0820_ ( .A1(\malu/Shift/_0069_ ), .A2(\malu/Shift/_0070_ ), .A3(\malu/Shift/_0717_ ), .ZN(\malu/Shift/_0071_ ) );
AOI21_X1 \malu/Shift/_0821_ ( .A(\malu/Shift/_0052_ ), .B1(\malu/Shift/_0067_ ), .B2(\malu/Shift/_0071_ ), .ZN(\malu/Shift/_0072_ ) );
AND2_X1 \malu/Shift/_0822_ ( .A1(\malu/Shift/_0042_ ), .A2(\malu/Shift/_0007_ ), .ZN(\malu/Shift/_0073_ ) );
AND2_X1 \malu/Shift/_0823_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0008_ ), .ZN(\malu/Shift/_0074_ ) );
OAI21_X1 \malu/Shift/_0824_ ( .A(\malu/Shift/_0033_ ), .B1(\malu/Shift/_0073_ ), .B2(\malu/Shift/_0074_ ), .ZN(\malu/Shift/_0075_ ) );
INV_X1 \malu/Shift/_0825_ ( .A(\malu/Shift/_0009_ ), .ZN(\malu/Shift/_0076_ ) );
NOR2_X1 \malu/Shift/_0826_ ( .A1(\malu/Shift/_0076_ ), .A2(\malu/Shift/_0716_ ), .ZN(\malu/Shift/_0077_ ) );
AND2_X1 \malu/Shift/_0827_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0010_ ), .ZN(\malu/Shift/_0078_ ) );
OAI21_X1 \malu/Shift/_0828_ ( .A(\malu/Shift/_0717_ ), .B1(\malu/Shift/_0077_ ), .B2(\malu/Shift/_0078_ ), .ZN(\malu/Shift/_0079_ ) );
BUF_X4 \malu/Shift/_0829_ ( .A(\malu/Shift/_0050_ ), .Z(\malu/Shift/_0080_ ) );
AND3_X1 \malu/Shift/_0830_ ( .A1(\malu/Shift/_0075_ ), .A2(\malu/Shift/_0079_ ), .A3(\malu/Shift/_0080_ ), .ZN(\malu/Shift/_0081_ ) );
OAI21_X1 \malu/Shift/_0831_ ( .A(\malu/Shift/_0064_ ), .B1(\malu/Shift/_0072_ ), .B2(\malu/Shift/_0081_ ), .ZN(\malu/Shift/_0082_ ) );
AND2_X4 \malu/Shift/_0832_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0017_ ), .ZN(\malu/Shift/_0083_ ) );
INV_X1 \malu/Shift/_0833_ ( .A(\malu/Shift/_0083_ ), .ZN(\malu/Shift/_0084_ ) );
INV_X1 \malu/Shift/_0834_ ( .A(\malu/Shift/_0016_ ), .ZN(\malu/Shift/_0085_ ) );
OAI211_X2 \malu/Shift/_0835_ ( .A(\malu/Shift/_0084_ ), .B(\malu/Shift/_0033_ ), .C1(\malu/Shift/_0716_ ), .C2(\malu/Shift/_0085_ ), .ZN(\malu/Shift/_0086_ ) );
AND2_X1 \malu/Shift/_0836_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0019_ ), .ZN(\malu/Shift/_0087_ ) );
INV_X1 \malu/Shift/_0837_ ( .A(\malu/Shift/_0087_ ), .ZN(\malu/Shift/_0088_ ) );
INV_X16 \malu/Shift/_0838_ ( .A(\malu/Shift/_0018_ ), .ZN(\malu/Shift/_0089_ ) );
OAI211_X2 \malu/Shift/_0839_ ( .A(\malu/Shift/_0088_ ), .B(\malu/Shift/_0717_ ), .C1(\malu/Shift/_0716_ ), .C2(\malu/Shift/_0089_ ), .ZN(\malu/Shift/_0090_ ) );
NAND3_X1 \malu/Shift/_0840_ ( .A1(\malu/Shift/_0086_ ), .A2(\malu/Shift/_0090_ ), .A3(\malu/Shift/_0080_ ), .ZN(\malu/Shift/_0091_ ) );
INV_X1 \malu/Shift/_0841_ ( .A(\malu/Shift/_0020_ ), .ZN(\malu/Shift/_0092_ ) );
NOR2_X1 \malu/Shift/_0842_ ( .A1(\malu/Shift/_0092_ ), .A2(\malu/Shift/_0716_ ), .ZN(\malu/Shift/_0093_ ) );
AND2_X1 \malu/Shift/_0843_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0021_ ), .ZN(\malu/Shift/_0094_ ) );
NOR2_X1 \malu/Shift/_0844_ ( .A1(\malu/Shift/_0093_ ), .A2(\malu/Shift/_0094_ ), .ZN(\malu/Shift/_0095_ ) );
INV_X16 \malu/Shift/_0845_ ( .A(\malu/Shift/_0023_ ), .ZN(\malu/Shift/_0096_ ) );
INV_X2 \malu/Shift/_0846_ ( .A(\malu/Shift/_0024_ ), .ZN(\malu/Shift/_0097_ ) );
MUX2_X1 \malu/Shift/_0847_ ( .A(\malu/Shift/_0096_ ), .B(\malu/Shift/_0097_ ), .S(\malu/Shift/_0716_ ), .Z(\malu/Shift/_0098_ ) );
MUX2_X1 \malu/Shift/_0848_ ( .A(\malu/Shift/_0095_ ), .B(\malu/Shift/_0098_ ), .S(\malu/Shift/_0717_ ), .Z(\malu/Shift/_0099_ ) );
BUF_X4 \malu/Shift/_0849_ ( .A(\malu/Shift/_0080_ ), .Z(\malu/Shift/_0100_ ) );
OAI211_X2 \malu/Shift/_0850_ ( .A(\malu/Shift/_0719_ ), .B(\malu/Shift/_0091_ ), .C1(\malu/Shift/_0099_ ), .C2(\malu/Shift/_0100_ ), .ZN(\malu/Shift/_0101_ ) );
AND3_X1 \malu/Shift/_0851_ ( .A1(\malu/Shift/_0082_ ), .A2(\malu/Shift/_0101_ ), .A3(\malu/Shift/_0720_ ), .ZN(\malu/Shift/_0102_ ) );
OAI21_X1 \malu/Shift/_0852_ ( .A(\malu/Shift/_0656_ ), .B1(\malu/Shift/_0063_ ), .B2(\malu/Shift/_0102_ ), .ZN(\malu/Shift/_0103_ ) );
INV_X1 \malu/Shift/_0853_ ( .A(\malu/Shift/_0635_ ), .ZN(\malu/Shift/_0104_ ) );
BUF_X4 \malu/Shift/_0854_ ( .A(\malu/Shift/_0104_ ), .Z(\malu/Shift/_0105_ ) );
AND3_X1 \malu/Shift/_0855_ ( .A1(\malu/Shift/_0032_ ), .A2(\malu/Shift/_0080_ ), .A3(\malu/Shift/_0039_ ), .ZN(\malu/Shift/_0106_ ) );
NAND2_X1 \malu/Shift/_0856_ ( .A1(\malu/Shift/_0106_ ), .A2(\malu/Shift/_0048_ ), .ZN(\malu/Shift/_0107_ ) );
INV_X1 \malu/Shift/_0857_ ( .A(\malu/Shift/_0720_ ), .ZN(\malu/Shift/_0108_ ) );
AND2_X1 \malu/Shift/_0858_ ( .A1(\malu/Shift/_0646_ ), .A2(\malu/Shift/_0108_ ), .ZN(\malu/Shift/_0109_ ) );
INV_X1 \malu/Shift/_0859_ ( .A(\malu/Shift/_0109_ ), .ZN(\malu/Shift/_0110_ ) );
OAI221_X1 \malu/Shift/_0860_ ( .A(\malu/Shift/_0103_ ), .B1(\malu/Shift/_0713_ ), .B2(\malu/Shift/_0105_ ), .C1(\malu/Shift/_0107_ ), .C2(\malu/Shift/_0110_ ), .ZN(\malu/Shift/_0721_ ) );
INV_X1 \malu/Shift/_0861_ ( .A(\malu/Shift/_0714_ ), .ZN(\malu/Shift/_0111_ ) );
NOR2_X1 \malu/Shift/_0862_ ( .A1(\malu/Shift/_0111_ ), .A2(\malu/Shift/_0715_ ), .ZN(\malu/Shift/_0112_ ) );
BUF_X4 \malu/Shift/_0863_ ( .A(\malu/Shift/_0112_ ), .Z(\malu/Shift/_0113_ ) );
AND2_X2 \malu/Shift/_0864_ ( .A1(\malu/Shift/_0042_ ), .A2(\malu/Shift/_0010_ ), .ZN(\malu/Shift/_0114_ ) );
INV_X1 \malu/Shift/_0865_ ( .A(\malu/Shift/_0114_ ), .ZN(\malu/Shift/_0115_ ) );
AND2_X1 \malu/Shift/_0866_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0012_ ), .ZN(\malu/Shift/_0116_ ) );
INV_X1 \malu/Shift/_0867_ ( .A(\malu/Shift/_0116_ ), .ZN(\malu/Shift/_0117_ ) );
NAND3_X1 \malu/Shift/_0868_ ( .A1(\malu/Shift/_0115_ ), .A2(\malu/Shift/_0717_ ), .A3(\malu/Shift/_0117_ ), .ZN(\malu/Shift/_0118_ ) );
AND2_X4 \malu/Shift/_0869_ ( .A1(\malu/Shift/_0042_ ), .A2(\malu/Shift/_0008_ ), .ZN(\malu/Shift/_0119_ ) );
INV_X1 \malu/Shift/_0870_ ( .A(\malu/Shift/_0119_ ), .ZN(\malu/Shift/_0120_ ) );
AND2_X1 \malu/Shift/_0871_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0009_ ), .ZN(\malu/Shift/_0121_ ) );
INV_X1 \malu/Shift/_0872_ ( .A(\malu/Shift/_0121_ ), .ZN(\malu/Shift/_0122_ ) );
NAND3_X1 \malu/Shift/_0873_ ( .A1(\malu/Shift/_0120_ ), .A2(\malu/Shift/_0033_ ), .A3(\malu/Shift/_0122_ ), .ZN(\malu/Shift/_0123_ ) );
AND3_X1 \malu/Shift/_0874_ ( .A1(\malu/Shift/_0118_ ), .A2(\malu/Shift/_0123_ ), .A3(\malu/Shift/_0050_ ), .ZN(\malu/Shift/_0124_ ) );
AND2_X2 \malu/Shift/_0875_ ( .A1(\malu/Shift/_0042_ ), .A2(\malu/Shift/_0013_ ), .ZN(\malu/Shift/_0125_ ) );
AND2_X1 \malu/Shift/_0876_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0014_ ), .ZN(\malu/Shift/_0126_ ) );
OAI21_X1 \malu/Shift/_0877_ ( .A(\malu/Shift/_0693_ ), .B1(\malu/Shift/_0125_ ), .B2(\malu/Shift/_0126_ ), .ZN(\malu/Shift/_0127_ ) );
AND2_X4 \malu/Shift/_0878_ ( .A1(\malu/Shift/_0042_ ), .A2(\malu/Shift/_0015_ ), .ZN(\malu/Shift/_0128_ ) );
AND2_X1 \malu/Shift/_0879_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0016_ ), .ZN(\malu/Shift/_0129_ ) );
OAI21_X1 \malu/Shift/_0880_ ( .A(\malu/Shift/_0717_ ), .B1(\malu/Shift/_0128_ ), .B2(\malu/Shift/_0129_ ), .ZN(\malu/Shift/_0130_ ) );
AOI21_X1 \malu/Shift/_0881_ ( .A(\malu/Shift/_0051_ ), .B1(\malu/Shift/_0127_ ), .B2(\malu/Shift/_0130_ ), .ZN(\malu/Shift/_0131_ ) );
NOR2_X1 \malu/Shift/_0882_ ( .A1(\malu/Shift/_0124_ ), .A2(\malu/Shift/_0131_ ), .ZN(\malu/Shift/_0132_ ) );
NOR2_X1 \malu/Shift/_0883_ ( .A1(\malu/Shift/_0132_ ), .A2(\malu/Shift/_0719_ ), .ZN(\malu/Shift/_0133_ ) );
INV_X1 \malu/Shift/_0884_ ( .A(\malu/Shift/_0021_ ), .ZN(\malu/Shift/_0134_ ) );
MUX2_X1 \malu/Shift/_0885_ ( .A(\malu/Shift/_0134_ ), .B(\malu/Shift/_0096_ ), .S(\malu/Shift/_0716_ ), .Z(\malu/Shift/_0135_ ) );
NOR2_X1 \malu/Shift/_0886_ ( .A1(\malu/Shift/_0135_ ), .A2(\malu/Shift/_0717_ ), .ZN(\malu/Shift/_0136_ ) );
AND2_X1 \malu/Shift/_0887_ ( .A1(\malu/Shift/_0717_ ), .A2(\malu/Shift/_0024_ ), .ZN(\malu/Shift/_0137_ ) );
OAI21_X1 \malu/Shift/_0888_ ( .A(\malu/Shift/_0718_ ), .B1(\malu/Shift/_0136_ ), .B2(\malu/Shift/_0137_ ), .ZN(\malu/Shift/_0138_ ) );
AND2_X2 \malu/Shift/_0889_ ( .A1(\malu/Shift/_0041_ ), .A2(\malu/Shift/_0017_ ), .ZN(\malu/Shift/_0139_ ) );
AND2_X1 \malu/Shift/_0890_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0018_ ), .ZN(\malu/Shift/_0140_ ) );
NOR2_X1 \malu/Shift/_0891_ ( .A1(\malu/Shift/_0139_ ), .A2(\malu/Shift/_0140_ ), .ZN(\malu/Shift/_0141_ ) );
AND2_X1 \malu/Shift/_0892_ ( .A1(\malu/Shift/_0041_ ), .A2(\malu/Shift/_0019_ ), .ZN(\malu/Shift/_0142_ ) );
AND2_X1 \malu/Shift/_0893_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0020_ ), .ZN(\malu/Shift/_0143_ ) );
NOR2_X2 \malu/Shift/_0894_ ( .A1(\malu/Shift/_0142_ ), .A2(\malu/Shift/_0143_ ), .ZN(\malu/Shift/_0144_ ) );
MUX2_X2 \malu/Shift/_0895_ ( .A(\malu/Shift/_0141_ ), .B(\malu/Shift/_0144_ ), .S(\malu/Shift/_0717_ ), .Z(\malu/Shift/_0145_ ) );
OAI21_X1 \malu/Shift/_0896_ ( .A(\malu/Shift/_0138_ ), .B1(\malu/Shift/_0145_ ), .B2(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0146_ ) );
AOI21_X1 \malu/Shift/_0897_ ( .A(\malu/Shift/_0133_ ), .B1(\malu/Shift/_0146_ ), .B2(\malu/Shift/_0719_ ), .ZN(\malu/Shift/_0147_ ) );
BUF_X2 \malu/Shift/_0898_ ( .A(\malu/Shift/_0108_ ), .Z(\malu/Shift/_0148_ ) );
BUF_X4 \malu/Shift/_0899_ ( .A(\malu/Shift/_0148_ ), .Z(\malu/Shift/_0149_ ) );
NOR2_X1 \malu/Shift/_0900_ ( .A1(\malu/Shift/_0147_ ), .A2(\malu/Shift/_0149_ ), .ZN(\malu/Shift/_0150_ ) );
BUF_X4 \malu/Shift/_0901_ ( .A(\malu/Shift/_0080_ ), .Z(\malu/Shift/_0151_ ) );
INV_X1 \malu/Shift/_0902_ ( .A(\malu/Shift/_0011_ ), .ZN(\malu/Shift/_0152_ ) );
NOR2_X1 \malu/Shift/_0903_ ( .A1(\malu/Shift/_0152_ ), .A2(\malu/Shift/_0716_ ), .ZN(\malu/Shift/_0153_ ) );
AND2_X1 \malu/Shift/_0904_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0022_ ), .ZN(\malu/Shift/_0154_ ) );
OR3_X1 \malu/Shift/_0905_ ( .A1(\malu/Shift/_0153_ ), .A2(\malu/Shift/_0154_ ), .A3(\malu/Shift/_0717_ ), .ZN(\malu/Shift/_0155_ ) );
AND2_X4 \malu/Shift/_0906_ ( .A1(\malu/Shift/_0042_ ), .A2(\malu/Shift/_0025_ ), .ZN(\malu/Shift/_0156_ ) );
AND2_X1 \malu/Shift/_0907_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0026_ ), .ZN(\malu/Shift/_0157_ ) );
NOR2_X1 \malu/Shift/_0908_ ( .A1(\malu/Shift/_0156_ ), .A2(\malu/Shift/_0157_ ), .ZN(\malu/Shift/_0158_ ) );
INV_X1 \malu/Shift/_0909_ ( .A(\malu/Shift/_0158_ ), .ZN(\malu/Shift/_0159_ ) );
OAI211_X2 \malu/Shift/_0910_ ( .A(\malu/Shift/_0151_ ), .B(\malu/Shift/_0155_ ), .C1(\malu/Shift/_0159_ ), .C2(\malu/Shift/_0039_ ), .ZN(\malu/Shift/_0160_ ) );
AND2_X2 \malu/Shift/_0911_ ( .A1(\malu/Shift/_0041_ ), .A2(\malu/Shift/_0029_ ), .ZN(\malu/Shift/_0161_ ) );
AND2_X4 \malu/Shift/_0912_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0030_ ), .ZN(\malu/Shift/_0162_ ) );
OR3_X1 \malu/Shift/_0913_ ( .A1(\malu/Shift/_0161_ ), .A2(\malu/Shift/_0034_ ), .A3(\malu/Shift/_0162_ ), .ZN(\malu/Shift/_0163_ ) );
AND2_X1 \malu/Shift/_0914_ ( .A1(\malu/Shift/_0042_ ), .A2(\malu/Shift/_0027_ ), .ZN(\malu/Shift/_0164_ ) );
INV_X1 \malu/Shift/_0915_ ( .A(\malu/Shift/_0164_ ), .ZN(\malu/Shift/_0165_ ) );
AND2_X4 \malu/Shift/_0916_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0028_ ), .ZN(\malu/Shift/_0166_ ) );
INV_X1 \malu/Shift/_0917_ ( .A(\malu/Shift/_0166_ ), .ZN(\malu/Shift/_0167_ ) );
NAND3_X1 \malu/Shift/_0918_ ( .A1(\malu/Shift/_0165_ ), .A2(\malu/Shift/_0039_ ), .A3(\malu/Shift/_0167_ ), .ZN(\malu/Shift/_0168_ ) );
NAND3_X1 \malu/Shift/_0919_ ( .A1(\malu/Shift/_0163_ ), .A2(\malu/Shift/_0168_ ), .A3(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0169_ ) );
NAND3_X1 \malu/Shift/_0920_ ( .A1(\malu/Shift/_0160_ ), .A2(\malu/Shift/_0064_ ), .A3(\malu/Shift/_0169_ ), .ZN(\malu/Shift/_0170_ ) );
INV_X1 \malu/Shift/_0921_ ( .A(\malu/Shift/_0004_ ), .ZN(\malu/Shift/_0171_ ) );
NOR2_X1 \malu/Shift/_0922_ ( .A1(\malu/Shift/_0171_ ), .A2(\malu/Shift/_0716_ ), .ZN(\malu/Shift/_0172_ ) );
AND2_X1 \malu/Shift/_0923_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0005_ ), .ZN(\malu/Shift/_0173_ ) );
OR3_X1 \malu/Shift/_0924_ ( .A1(\malu/Shift/_0172_ ), .A2(\malu/Shift/_0173_ ), .A3(\malu/Shift/_0717_ ), .ZN(\malu/Shift/_0174_ ) );
INV_X1 \malu/Shift/_0925_ ( .A(\malu/Shift/_0006_ ), .ZN(\malu/Shift/_0175_ ) );
NOR2_X1 \malu/Shift/_0926_ ( .A1(\malu/Shift/_0175_ ), .A2(\malu/Shift/_0716_ ), .ZN(\malu/Shift/_0176_ ) );
INV_X1 \malu/Shift/_0927_ ( .A(\malu/Shift/_0176_ ), .ZN(\malu/Shift/_0177_ ) );
AND2_X1 \malu/Shift/_0928_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0007_ ), .ZN(\malu/Shift/_0178_ ) );
INV_X1 \malu/Shift/_0929_ ( .A(\malu/Shift/_0178_ ), .ZN(\malu/Shift/_0179_ ) );
NAND3_X1 \malu/Shift/_0930_ ( .A1(\malu/Shift/_0177_ ), .A2(\malu/Shift/_0717_ ), .A3(\malu/Shift/_0179_ ), .ZN(\malu/Shift/_0180_ ) );
AOI21_X1 \malu/Shift/_0931_ ( .A(\malu/Shift/_0080_ ), .B1(\malu/Shift/_0174_ ), .B2(\malu/Shift/_0180_ ), .ZN(\malu/Shift/_0181_ ) );
INV_X1 \malu/Shift/_0932_ ( .A(\malu/Shift/_0031_ ), .ZN(\malu/Shift/_0182_ ) );
NOR2_X1 \malu/Shift/_0933_ ( .A1(\malu/Shift/_0182_ ), .A2(\malu/Shift/_0716_ ), .ZN(\malu/Shift/_0183_ ) );
AND2_X1 \malu/Shift/_0934_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0001_ ), .ZN(\malu/Shift/_0184_ ) );
OAI21_X1 \malu/Shift/_0935_ ( .A(\malu/Shift/_0038_ ), .B1(\malu/Shift/_0183_ ), .B2(\malu/Shift/_0184_ ), .ZN(\malu/Shift/_0185_ ) );
INV_X1 \malu/Shift/_0936_ ( .A(\malu/Shift/_0002_ ), .ZN(\malu/Shift/_0186_ ) );
NOR2_X1 \malu/Shift/_0937_ ( .A1(\malu/Shift/_0186_ ), .A2(\malu/Shift/_0716_ ), .ZN(\malu/Shift/_0187_ ) );
AND2_X1 \malu/Shift/_0938_ ( .A1(\malu/Shift/_0716_ ), .A2(\malu/Shift/_0003_ ), .ZN(\malu/Shift/_0188_ ) );
OAI21_X1 \malu/Shift/_0939_ ( .A(\malu/Shift/_0717_ ), .B1(\malu/Shift/_0187_ ), .B2(\malu/Shift/_0188_ ), .ZN(\malu/Shift/_0189_ ) );
AND3_X1 \malu/Shift/_0940_ ( .A1(\malu/Shift/_0185_ ), .A2(\malu/Shift/_0189_ ), .A3(\malu/Shift/_0051_ ), .ZN(\malu/Shift/_0190_ ) );
OAI21_X1 \malu/Shift/_0941_ ( .A(\malu/Shift/_0719_ ), .B1(\malu/Shift/_0181_ ), .B2(\malu/Shift/_0190_ ), .ZN(\malu/Shift/_0191_ ) );
AND3_X1 \malu/Shift/_0942_ ( .A1(\malu/Shift/_0170_ ), .A2(\malu/Shift/_0191_ ), .A3(\malu/Shift/_0148_ ), .ZN(\malu/Shift/_0192_ ) );
OAI21_X1 \malu/Shift/_0943_ ( .A(\malu/Shift/_0113_ ), .B1(\malu/Shift/_0150_ ), .B2(\malu/Shift/_0192_ ), .ZN(\malu/Shift/_0193_ ) );
AND2_X2 \malu/Shift/_0944_ ( .A1(\malu/Shift/_0111_ ), .A2(\malu/Shift/_0715_ ), .ZN(\malu/Shift/_0194_ ) );
NAND4_X1 \malu/Shift/_0945_ ( .A1(\malu/Shift/_0170_ ), .A2(\malu/Shift/_0191_ ), .A3(\malu/Shift/_0149_ ), .A4(\malu/Shift/_0194_ ), .ZN(\malu/Shift/_0195_ ) );
AND2_X1 \malu/Shift/_0946_ ( .A1(\malu/Shift/_0194_ ), .A2(\malu/Shift/_0720_ ), .ZN(\malu/Shift/_0196_ ) );
NOR2_X1 \malu/Shift/_0947_ ( .A1(\malu/Shift/_0097_ ), .A2(\malu/Shift/_0716_ ), .ZN(\malu/Shift/_0197_ ) );
AOI21_X1 \malu/Shift/_0948_ ( .A(\malu/Shift/_0136_ ), .B1(\malu/Shift/_0717_ ), .B2(\malu/Shift/_0197_ ), .ZN(\malu/Shift/_0198_ ) );
MUX2_X1 \malu/Shift/_0949_ ( .A(\malu/Shift/_0145_ ), .B(\malu/Shift/_0198_ ), .S(\malu/Shift/_0718_ ), .Z(\malu/Shift/_0199_ ) );
NOR2_X1 \malu/Shift/_0950_ ( .A1(\malu/Shift/_0199_ ), .A2(\malu/Shift/_0048_ ), .ZN(\malu/Shift/_0200_ ) );
OAI21_X1 \malu/Shift/_0951_ ( .A(\malu/Shift/_0196_ ), .B1(\malu/Shift/_0200_ ), .B2(\malu/Shift/_0133_ ), .ZN(\malu/Shift/_0201_ ) );
MUX2_X1 \malu/Shift/_0952_ ( .A(\malu/Shift/_0152_ ), .B(\malu/Shift/_0713_ ), .S(\malu/Shift/_0716_ ), .Z(\malu/Shift/_0202_ ) );
NOR3_X1 \malu/Shift/_0953_ ( .A1(\malu/Shift/_0202_ ), .A2(\malu/Shift/_0718_ ), .A3(\malu/Shift/_0717_ ), .ZN(\malu/Shift/_0203_ ) );
AND2_X1 \malu/Shift/_0954_ ( .A1(\malu/Shift/_0203_ ), .A2(\malu/Shift/_0064_ ), .ZN(\malu/Shift/_0204_ ) );
BUF_X2 \malu/Shift/_0955_ ( .A(\malu/Shift/_0109_ ), .Z(\malu/Shift/_0205_ ) );
AOI22_X1 \malu/Shift/_0956_ ( .A1(\malu/Shift/_0204_ ), .A2(\malu/Shift/_0205_ ), .B1(\malu/Shift/_0011_ ), .B2(\malu/Shift/_0635_ ), .ZN(\malu/Shift/_0206_ ) );
NAND4_X1 \malu/Shift/_0957_ ( .A1(\malu/Shift/_0193_ ), .A2(\malu/Shift/_0195_ ), .A3(\malu/Shift/_0201_ ), .A4(\malu/Shift/_0206_ ), .ZN(\malu/Shift/_0732_ ) );
OR3_X4 \malu/Shift/_0958_ ( .A1(\malu/Shift/_0069_ ), .A2(\malu/Shift/_0070_ ), .A3(\malu/Shift/_0693_ ), .ZN(\malu/Shift/_0207_ ) );
INV_X1 \malu/Shift/_0959_ ( .A(\malu/Shift/_0078_ ), .ZN(\malu/Shift/_0208_ ) );
OAI211_X2 \malu/Shift/_0960_ ( .A(\malu/Shift/_0208_ ), .B(\malu/Shift/_0693_ ), .C1(\malu/Shift/_0716_ ), .C2(\malu/Shift/_0076_ ), .ZN(\malu/Shift/_0209_ ) );
NAND3_X1 \malu/Shift/_0961_ ( .A1(\malu/Shift/_0207_ ), .A2(\malu/Shift/_0209_ ), .A3(\malu/Shift/_0050_ ), .ZN(\malu/Shift/_0210_ ) );
OR3_X2 \malu/Shift/_0962_ ( .A1(\malu/Shift/_0065_ ), .A2(\malu/Shift/_0066_ ), .A3(\malu/Shift/_0717_ ), .ZN(\malu/Shift/_0211_ ) );
OAI211_X2 \malu/Shift/_0963_ ( .A(\malu/Shift/_0084_ ), .B(\malu/Shift/_0717_ ), .C1(\malu/Shift/_0716_ ), .C2(\malu/Shift/_0085_ ), .ZN(\malu/Shift/_0212_ ) );
AND2_X2 \malu/Shift/_0964_ ( .A1(\malu/Shift/_0211_ ), .A2(\malu/Shift/_0212_ ), .ZN(\malu/Shift/_0213_ ) );
INV_X2 \malu/Shift/_0965_ ( .A(\malu/Shift/_0213_ ), .ZN(\malu/Shift/_0214_ ) );
OAI21_X1 \malu/Shift/_0966_ ( .A(\malu/Shift/_0210_ ), .B1(\malu/Shift/_0214_ ), .B2(\malu/Shift/_0050_ ), .ZN(\malu/Shift/_0215_ ) );
AND2_X2 \malu/Shift/_0967_ ( .A1(\malu/Shift/_0215_ ), .A2(\malu/Shift/_0710_ ), .ZN(\malu/Shift/_0216_ ) );
NOR2_X1 \malu/Shift/_0968_ ( .A1(\malu/Shift/_0089_ ), .A2(\malu/Shift/_0716_ ), .ZN(\malu/Shift/_0217_ ) );
NOR2_X1 \malu/Shift/_0969_ ( .A1(\malu/Shift/_0217_ ), .A2(\malu/Shift/_0087_ ), .ZN(\malu/Shift/_0218_ ) );
MUX2_X1 \malu/Shift/_0970_ ( .A(\malu/Shift/_0218_ ), .B(\malu/Shift/_0095_ ), .S(\malu/Shift/_0717_ ), .Z(\malu/Shift/_0219_ ) );
OR2_X1 \malu/Shift/_0971_ ( .A1(\malu/Shift/_0219_ ), .A2(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0220_ ) );
NAND3_X1 \malu/Shift/_0972_ ( .A1(\malu/Shift/_0718_ ), .A2(\malu/Shift/_0717_ ), .A3(\malu/Shift/_0024_ ), .ZN(\malu/Shift/_0221_ ) );
OR3_X1 \malu/Shift/_0973_ ( .A1(\malu/Shift/_0098_ ), .A2(\malu/Shift/_0050_ ), .A3(\malu/Shift/_0717_ ), .ZN(\malu/Shift/_0222_ ) );
NAND3_X2 \malu/Shift/_0974_ ( .A1(\malu/Shift/_0220_ ), .A2(\malu/Shift/_0221_ ), .A3(\malu/Shift/_0222_ ), .ZN(\malu/Shift/_0223_ ) );
AOI21_X2 \malu/Shift/_0975_ ( .A(\malu/Shift/_0216_ ), .B1(\malu/Shift/_0223_ ), .B2(\malu/Shift/_0719_ ), .ZN(\malu/Shift/_0224_ ) );
NOR2_X1 \malu/Shift/_0976_ ( .A1(\malu/Shift/_0224_ ), .A2(\malu/Shift/_0148_ ), .ZN(\malu/Shift/_0225_ ) );
OR3_X1 \malu/Shift/_0977_ ( .A1(\malu/Shift/_0702_ ), .A2(\malu/Shift/_0703_ ), .A3(\malu/Shift/_0700_ ), .ZN(\malu/Shift/_0226_ ) );
OR3_X1 \malu/Shift/_0978_ ( .A1(\malu/Shift/_0676_ ), .A2(\malu/Shift/_0686_ ), .A3(\malu/Shift/_0717_ ), .ZN(\malu/Shift/_0227_ ) );
AOI21_X1 \malu/Shift/_0979_ ( .A(\malu/Shift/_0718_ ), .B1(\malu/Shift/_0226_ ), .B2(\malu/Shift/_0227_ ), .ZN(\malu/Shift/_0228_ ) );
OAI21_X1 \malu/Shift/_0980_ ( .A(\malu/Shift/_0717_ ), .B1(\malu/Shift/_0073_ ), .B2(\malu/Shift/_0074_ ), .ZN(\malu/Shift/_0229_ ) );
OAI21_X1 \malu/Shift/_0981_ ( .A(\malu/Shift/_0700_ ), .B1(\malu/Shift/_0706_ ), .B2(\malu/Shift/_0707_ ), .ZN(\malu/Shift/_0230_ ) );
AND3_X1 \malu/Shift/_0982_ ( .A1(\malu/Shift/_0229_ ), .A2(\malu/Shift/_0718_ ), .A3(\malu/Shift/_0230_ ), .ZN(\malu/Shift/_0231_ ) );
NOR2_X1 \malu/Shift/_0983_ ( .A1(\malu/Shift/_0228_ ), .A2(\malu/Shift/_0231_ ), .ZN(\malu/Shift/_0232_ ) );
NAND2_X1 \malu/Shift/_0984_ ( .A1(\malu/Shift/_0232_ ), .A2(\malu/Shift/_0719_ ), .ZN(\malu/Shift/_0233_ ) );
OAI21_X1 \malu/Shift/_0985_ ( .A(\malu/Shift/_0717_ ), .B1(\malu/Shift/_0054_ ), .B2(\malu/Shift/_0055_ ), .ZN(\malu/Shift/_0234_ ) );
OAI211_X2 \malu/Shift/_0986_ ( .A(\malu/Shift/_0234_ ), .B(\malu/Shift/_0100_ ), .C1(\malu/Shift/_0045_ ), .C2(\malu/Shift/_0717_ ), .ZN(\malu/Shift/_0235_ ) );
BUF_X4 \malu/Shift/_0987_ ( .A(\malu/Shift/_0047_ ), .Z(\malu/Shift/_0236_ ) );
OAI21_X1 \malu/Shift/_0988_ ( .A(\malu/Shift/_0038_ ), .B1(\malu/Shift/_0058_ ), .B2(\malu/Shift/_0059_ ), .ZN(\malu/Shift/_0237_ ) );
OAI21_X1 \malu/Shift/_0989_ ( .A(\malu/Shift/_0717_ ), .B1(\malu/Shift/_0696_ ), .B2(\malu/Shift/_0697_ ), .ZN(\malu/Shift/_0238_ ) );
NAND2_X1 \malu/Shift/_0990_ ( .A1(\malu/Shift/_0237_ ), .A2(\malu/Shift/_0238_ ), .ZN(\malu/Shift/_0239_ ) );
OAI211_X2 \malu/Shift/_0991_ ( .A(\malu/Shift/_0235_ ), .B(\malu/Shift/_0236_ ), .C1(\malu/Shift/_0053_ ), .C2(\malu/Shift/_0239_ ), .ZN(\malu/Shift/_0240_ ) );
AOI21_X1 \malu/Shift/_0992_ ( .A(\malu/Shift/_0720_ ), .B1(\malu/Shift/_0233_ ), .B2(\malu/Shift/_0240_ ), .ZN(\malu/Shift/_0241_ ) );
OAI21_X1 \malu/Shift/_0993_ ( .A(\malu/Shift/_0113_ ), .B1(\malu/Shift/_0225_ ), .B2(\malu/Shift/_0241_ ), .ZN(\malu/Shift/_0242_ ) );
NAND2_X1 \malu/Shift/_0994_ ( .A1(\malu/Shift/_0241_ ), .A2(\malu/Shift/_0194_ ), .ZN(\malu/Shift/_0243_ ) );
AOI21_X1 \malu/Shift/_0995_ ( .A(\malu/Shift/_0711_ ), .B1(\malu/Shift/_0220_ ), .B2(\malu/Shift/_0222_ ), .ZN(\malu/Shift/_0244_ ) );
OAI21_X1 \malu/Shift/_0996_ ( .A(\malu/Shift/_0196_ ), .B1(\malu/Shift/_0216_ ), .B2(\malu/Shift/_0244_ ), .ZN(\malu/Shift/_0245_ ) );
OR3_X4 \malu/Shift/_0997_ ( .A1(\malu/Shift/_0043_ ), .A2(\malu/Shift/_0037_ ), .A3(\malu/Shift/_0717_ ), .ZN(\malu/Shift/_0246_ ) );
OAI21_X2 \malu/Shift/_0998_ ( .A(\malu/Shift/_0246_ ), .B1(\malu/Shift/_0033_ ), .B2(\malu/Shift/_0032_ ), .ZN(\malu/Shift/_0247_ ) );
NOR4_X1 \malu/Shift/_0999_ ( .A1(\malu/Shift/_0247_ ), .A2(\malu/Shift/_0720_ ), .A3(\malu/Shift/_0718_ ), .A4(\malu/Shift/_0719_ ), .ZN(\malu/Shift/_0248_ ) );
BUF_X2 \malu/Shift/_1000_ ( .A(\malu/Shift/_0646_ ), .Z(\malu/Shift/_0249_ ) );
AOI22_X1 \malu/Shift/_1001_ ( .A1(\malu/Shift/_0248_ ), .A2(\malu/Shift/_0249_ ), .B1(\malu/Shift/_0022_ ), .B2(\malu/Shift/_0635_ ), .ZN(\malu/Shift/_0250_ ) );
NAND4_X1 \malu/Shift/_1002_ ( .A1(\malu/Shift/_0242_ ), .A2(\malu/Shift/_0243_ ), .A3(\malu/Shift/_0245_ ), .A4(\malu/Shift/_0250_ ), .ZN(\malu/Shift/_0743_ ) );
MUX2_X1 \malu/Shift/_1003_ ( .A(\malu/Shift/_0135_ ), .B(\malu/Shift/_0144_ ), .S(\malu/Shift/_0700_ ), .Z(\malu/Shift/_0251_ ) );
OR2_X2 \malu/Shift/_1004_ ( .A1(\malu/Shift/_0251_ ), .A2(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0252_ ) );
AND2_X1 \malu/Shift/_1005_ ( .A1(\malu/Shift/_0718_ ), .A2(\malu/Shift/_0024_ ), .ZN(\malu/Shift/_0253_ ) );
INV_X1 \malu/Shift/_1006_ ( .A(\malu/Shift/_0253_ ), .ZN(\malu/Shift/_0254_ ) );
AOI21_X1 \malu/Shift/_1007_ ( .A(\malu/Shift/_0064_ ), .B1(\malu/Shift/_0252_ ), .B2(\malu/Shift/_0254_ ), .ZN(\malu/Shift/_0255_ ) );
OR3_X1 \malu/Shift/_1008_ ( .A1(\malu/Shift/_0139_ ), .A2(\malu/Shift/_0700_ ), .A3(\malu/Shift/_0140_ ), .ZN(\malu/Shift/_0256_ ) );
OR3_X1 \malu/Shift/_1009_ ( .A1(\malu/Shift/_0128_ ), .A2(\malu/Shift/_0717_ ), .A3(\malu/Shift/_0129_ ), .ZN(\malu/Shift/_0257_ ) );
NAND3_X1 \malu/Shift/_1010_ ( .A1(\malu/Shift/_0256_ ), .A2(\malu/Shift/_0257_ ), .A3(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0258_ ) );
OR3_X1 \malu/Shift/_1011_ ( .A1(\malu/Shift/_0125_ ), .A2(\malu/Shift/_0700_ ), .A3(\malu/Shift/_0126_ ), .ZN(\malu/Shift/_0259_ ) );
NAND3_X1 \malu/Shift/_1012_ ( .A1(\malu/Shift/_0115_ ), .A2(\malu/Shift/_0033_ ), .A3(\malu/Shift/_0117_ ), .ZN(\malu/Shift/_0260_ ) );
NAND3_X1 \malu/Shift/_1013_ ( .A1(\malu/Shift/_0259_ ), .A2(\malu/Shift/_0260_ ), .A3(\malu/Shift/_0051_ ), .ZN(\malu/Shift/_0261_ ) );
AOI21_X1 \malu/Shift/_1014_ ( .A(\malu/Shift/_0719_ ), .B1(\malu/Shift/_0258_ ), .B2(\malu/Shift/_0261_ ), .ZN(\malu/Shift/_0262_ ) );
NOR2_X1 \malu/Shift/_1015_ ( .A1(\malu/Shift/_0255_ ), .A2(\malu/Shift/_0262_ ), .ZN(\malu/Shift/_0263_ ) );
NOR2_X1 \malu/Shift/_1016_ ( .A1(\malu/Shift/_0263_ ), .A2(\malu/Shift/_0148_ ), .ZN(\malu/Shift/_0264_ ) );
NAND3_X1 \malu/Shift/_1017_ ( .A1(\malu/Shift/_0165_ ), .A2(\malu/Shift/_0717_ ), .A3(\malu/Shift/_0167_ ), .ZN(\malu/Shift/_0265_ ) );
OAI211_X2 \malu/Shift/_1018_ ( .A(\malu/Shift/_0151_ ), .B(\malu/Shift/_0265_ ), .C1(\malu/Shift/_0159_ ), .C2(\malu/Shift/_0717_ ), .ZN(\malu/Shift/_0266_ ) );
OR3_X1 \malu/Shift/_1019_ ( .A1(\malu/Shift/_0161_ ), .A2(\malu/Shift/_0717_ ), .A3(\malu/Shift/_0162_ ), .ZN(\malu/Shift/_0267_ ) );
OR3_X1 \malu/Shift/_1020_ ( .A1(\malu/Shift/_0183_ ), .A2(\malu/Shift/_0184_ ), .A3(\malu/Shift/_0038_ ), .ZN(\malu/Shift/_0268_ ) );
NAND2_X1 \malu/Shift/_1021_ ( .A1(\malu/Shift/_0267_ ), .A2(\malu/Shift/_0268_ ), .ZN(\malu/Shift/_0269_ ) );
OAI211_X2 \malu/Shift/_1022_ ( .A(\malu/Shift/_0266_ ), .B(\malu/Shift/_0064_ ), .C1(\malu/Shift/_0269_ ), .C2(\malu/Shift/_0100_ ), .ZN(\malu/Shift/_0270_ ) );
OAI21_X1 \malu/Shift/_1023_ ( .A(\malu/Shift/_0038_ ), .B1(\malu/Shift/_0187_ ), .B2(\malu/Shift/_0188_ ), .ZN(\malu/Shift/_0271_ ) );
OAI21_X1 \malu/Shift/_1024_ ( .A(\malu/Shift/_0717_ ), .B1(\malu/Shift/_0172_ ), .B2(\malu/Shift/_0173_ ), .ZN(\malu/Shift/_0272_ ) );
NAND2_X1 \malu/Shift/_1025_ ( .A1(\malu/Shift/_0271_ ), .A2(\malu/Shift/_0272_ ), .ZN(\malu/Shift/_0273_ ) );
NAND2_X1 \malu/Shift/_1026_ ( .A1(\malu/Shift/_0273_ ), .A2(\malu/Shift/_0052_ ), .ZN(\malu/Shift/_0274_ ) );
NAND3_X1 \malu/Shift/_1027_ ( .A1(\malu/Shift/_0120_ ), .A2(\malu/Shift/_0717_ ), .A3(\malu/Shift/_0122_ ), .ZN(\malu/Shift/_0275_ ) );
NAND3_X1 \malu/Shift/_1028_ ( .A1(\malu/Shift/_0177_ ), .A2(\malu/Shift/_0034_ ), .A3(\malu/Shift/_0179_ ), .ZN(\malu/Shift/_0276_ ) );
NAND3_X1 \malu/Shift/_1029_ ( .A1(\malu/Shift/_0275_ ), .A2(\malu/Shift/_0718_ ), .A3(\malu/Shift/_0276_ ), .ZN(\malu/Shift/_0277_ ) );
NAND3_X1 \malu/Shift/_1030_ ( .A1(\malu/Shift/_0274_ ), .A2(\malu/Shift/_0277_ ), .A3(\malu/Shift/_0719_ ), .ZN(\malu/Shift/_0278_ ) );
AND3_X1 \malu/Shift/_1031_ ( .A1(\malu/Shift/_0270_ ), .A2(\malu/Shift/_0148_ ), .A3(\malu/Shift/_0278_ ), .ZN(\malu/Shift/_0279_ ) );
OAI21_X1 \malu/Shift/_1032_ ( .A(\malu/Shift/_0113_ ), .B1(\malu/Shift/_0264_ ), .B2(\malu/Shift/_0279_ ), .ZN(\malu/Shift/_0280_ ) );
NAND4_X1 \malu/Shift/_1033_ ( .A1(\malu/Shift/_0270_ ), .A2(\malu/Shift/_0149_ ), .A3(\malu/Shift/_0194_ ), .A4(\malu/Shift/_0278_ ), .ZN(\malu/Shift/_0281_ ) );
NOR3_X1 \malu/Shift/_1034_ ( .A1(\malu/Shift/_0097_ ), .A2(\malu/Shift/_0717_ ), .A3(\malu/Shift/_0716_ ), .ZN(\malu/Shift/_0282_ ) );
INV_X1 \malu/Shift/_1035_ ( .A(\malu/Shift/_0282_ ), .ZN(\malu/Shift/_0283_ ) );
OAI21_X1 \malu/Shift/_1036_ ( .A(\malu/Shift/_0252_ ), .B1(\malu/Shift/_0052_ ), .B2(\malu/Shift/_0283_ ), .ZN(\malu/Shift/_0284_ ) );
AND2_X1 \malu/Shift/_1037_ ( .A1(\malu/Shift/_0284_ ), .A2(\malu/Shift/_0719_ ), .ZN(\malu/Shift/_0285_ ) );
OAI21_X1 \malu/Shift/_1038_ ( .A(\malu/Shift/_0196_ ), .B1(\malu/Shift/_0285_ ), .B2(\malu/Shift/_0262_ ), .ZN(\malu/Shift/_0286_ ) );
NOR2_X1 \malu/Shift/_1039_ ( .A1(\malu/Shift/_0156_ ), .A2(\malu/Shift/_0154_ ), .ZN(\malu/Shift/_0287_ ) );
MUX2_X2 \malu/Shift/_1040_ ( .A(\malu/Shift/_0202_ ), .B(\malu/Shift/_0287_ ), .S(\malu/Shift/_0700_ ), .Z(\malu/Shift/_0288_ ) );
NOR2_X1 \malu/Shift/_1041_ ( .A1(\malu/Shift/_0288_ ), .A2(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0289_ ) );
AND2_X1 \malu/Shift/_1042_ ( .A1(\malu/Shift/_0289_ ), .A2(\malu/Shift/_0047_ ), .ZN(\malu/Shift/_0290_ ) );
AOI22_X1 \malu/Shift/_1043_ ( .A1(\malu/Shift/_0290_ ), .A2(\malu/Shift/_0205_ ), .B1(\malu/Shift/_0025_ ), .B2(\malu/Shift/_0635_ ), .ZN(\malu/Shift/_0291_ ) );
NAND4_X1 \malu/Shift/_1044_ ( .A1(\malu/Shift/_0280_ ), .A2(\malu/Shift/_0281_ ), .A3(\malu/Shift/_0286_ ), .A4(\malu/Shift/_0291_ ), .ZN(\malu/Shift/_0746_ ) );
NAND3_X1 \malu/Shift/_1045_ ( .A1(\malu/Shift/_0714_ ), .A2(\malu/Shift/_0715_ ), .A3(\malu/Shift/_0026_ ), .ZN(\malu/Shift/_0292_ ) );
OAI21_X1 \malu/Shift/_1046_ ( .A(\malu/Shift/_0700_ ), .B1(\malu/Shift/_0054_ ), .B2(\malu/Shift/_0044_ ), .ZN(\malu/Shift/_0293_ ) );
OAI21_X1 \malu/Shift/_1047_ ( .A(\malu/Shift/_0717_ ), .B1(\malu/Shift/_0043_ ), .B2(\malu/Shift/_0037_ ), .ZN(\malu/Shift/_0294_ ) );
NAND2_X1 \malu/Shift/_1048_ ( .A1(\malu/Shift/_0293_ ), .A2(\malu/Shift/_0294_ ), .ZN(\malu/Shift/_0295_ ) );
NAND2_X1 \malu/Shift/_1049_ ( .A1(\malu/Shift/_0295_ ), .A2(\malu/Shift/_0051_ ), .ZN(\malu/Shift/_0296_ ) );
NAND4_X1 \malu/Shift/_1050_ ( .A1(\malu/Shift/_0038_ ), .A2(\malu/Shift/_0042_ ), .A3(\malu/Shift/_0718_ ), .A4(\malu/Shift/_0000_ ), .ZN(\malu/Shift/_0297_ ) );
NAND2_X1 \malu/Shift/_1051_ ( .A1(\malu/Shift/_0296_ ), .A2(\malu/Shift/_0297_ ), .ZN(\malu/Shift/_0298_ ) );
AND3_X1 \malu/Shift/_1052_ ( .A1(\malu/Shift/_0298_ ), .A2(\malu/Shift/_0711_ ), .A3(\malu/Shift/_0646_ ), .ZN(\malu/Shift/_0299_ ) );
AOI21_X1 \malu/Shift/_1053_ ( .A(\malu/Shift/_0050_ ), .B1(\malu/Shift/_0075_ ), .B2(\malu/Shift/_0079_ ), .ZN(\malu/Shift/_0300_ ) );
AOI21_X1 \malu/Shift/_1054_ ( .A(\malu/Shift/_0718_ ), .B1(\malu/Shift/_0704_ ), .B2(\malu/Shift/_0708_ ), .ZN(\malu/Shift/_0301_ ) );
OR2_X1 \malu/Shift/_1055_ ( .A1(\malu/Shift/_0300_ ), .A2(\malu/Shift/_0301_ ), .ZN(\malu/Shift/_0302_ ) );
AND2_X2 \malu/Shift/_1056_ ( .A1(\malu/Shift/_0694_ ), .A2(\malu/Shift/_0698_ ), .ZN(\malu/Shift/_0303_ ) );
MUX2_X2 \malu/Shift/_1057_ ( .A(\malu/Shift/_0061_ ), .B(\malu/Shift/_0303_ ), .S(\malu/Shift/_0718_ ), .Z(\malu/Shift/_0304_ ) );
MUX2_X2 \malu/Shift/_1058_ ( .A(\malu/Shift/_0302_ ), .B(\malu/Shift/_0304_ ), .S(\malu/Shift/_0711_ ), .Z(\malu/Shift/_0305_ ) );
OR2_X2 \malu/Shift/_1059_ ( .A1(\malu/Shift/_0305_ ), .A2(\malu/Shift/_0720_ ), .ZN(\malu/Shift/_0306_ ) );
AOI21_X1 \malu/Shift/_1060_ ( .A(\malu/Shift/_0299_ ), .B1(\malu/Shift/_0306_ ), .B2(\malu/Shift/_0656_ ), .ZN(\malu/Shift/_0307_ ) );
INV_X1 \malu/Shift/_1061_ ( .A(\malu/Shift/_0112_ ), .ZN(\malu/Shift/_0308_ ) );
NOR2_X1 \malu/Shift/_1062_ ( .A1(\malu/Shift/_0099_ ), .A2(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0309_ ) );
OAI21_X1 \malu/Shift/_1063_ ( .A(\malu/Shift/_0719_ ), .B1(\malu/Shift/_0309_ ), .B2(\malu/Shift/_0253_ ), .ZN(\malu/Shift/_0310_ ) );
AOI21_X1 \malu/Shift/_1064_ ( .A(\malu/Shift/_0718_ ), .B1(\malu/Shift/_0067_ ), .B2(\malu/Shift/_0071_ ), .ZN(\malu/Shift/_0311_ ) );
AOI21_X1 \malu/Shift/_1065_ ( .A(\malu/Shift/_0050_ ), .B1(\malu/Shift/_0086_ ), .B2(\malu/Shift/_0090_ ), .ZN(\malu/Shift/_0312_ ) );
NOR2_X1 \malu/Shift/_1066_ ( .A1(\malu/Shift/_0311_ ), .A2(\malu/Shift/_0312_ ), .ZN(\malu/Shift/_0313_ ) );
NAND2_X1 \malu/Shift/_1067_ ( .A1(\malu/Shift/_0313_ ), .A2(\malu/Shift/_0236_ ), .ZN(\malu/Shift/_0314_ ) );
AOI21_X1 \malu/Shift/_1068_ ( .A(\malu/Shift/_0308_ ), .B1(\malu/Shift/_0310_ ), .B2(\malu/Shift/_0314_ ), .ZN(\malu/Shift/_0315_ ) );
INV_X1 \malu/Shift/_1069_ ( .A(\malu/Shift/_0194_ ), .ZN(\malu/Shift/_0316_ ) );
OR3_X1 \malu/Shift/_1070_ ( .A1(\malu/Shift/_0099_ ), .A2(\malu/Shift/_0718_ ), .A3(\malu/Shift/_0047_ ), .ZN(\malu/Shift/_0317_ ) );
AOI21_X1 \malu/Shift/_1071_ ( .A(\malu/Shift/_0316_ ), .B1(\malu/Shift/_0314_ ), .B2(\malu/Shift/_0317_ ), .ZN(\malu/Shift/_0318_ ) );
NOR3_X1 \malu/Shift/_1072_ ( .A1(\malu/Shift/_0315_ ), .A2(\malu/Shift/_0318_ ), .A3(\malu/Shift/_0149_ ), .ZN(\malu/Shift/_0319_ ) );
OAI21_X1 \malu/Shift/_1073_ ( .A(\malu/Shift/_0292_ ), .B1(\malu/Shift/_0307_ ), .B2(\malu/Shift/_0319_ ), .ZN(\malu/Shift/_0747_ ) );
OR3_X1 \malu/Shift/_1074_ ( .A1(\malu/Shift/_0198_ ), .A2(\malu/Shift/_0718_ ), .A3(\malu/Shift/_0710_ ), .ZN(\malu/Shift/_0320_ ) );
AND2_X1 \malu/Shift/_1075_ ( .A1(\malu/Shift/_0127_ ), .A2(\malu/Shift/_0130_ ), .ZN(\malu/Shift/_0321_ ) );
MUX2_X2 \malu/Shift/_1076_ ( .A(\malu/Shift/_0321_ ), .B(\malu/Shift/_0145_ ), .S(\malu/Shift/_0718_ ), .Z(\malu/Shift/_0322_ ) );
OAI21_X1 \malu/Shift/_1077_ ( .A(\malu/Shift/_0320_ ), .B1(\malu/Shift/_0322_ ), .B2(\malu/Shift/_0719_ ), .ZN(\malu/Shift/_0323_ ) );
NAND2_X1 \malu/Shift/_1078_ ( .A1(\malu/Shift/_0323_ ), .A2(\malu/Shift/_0194_ ), .ZN(\malu/Shift/_0324_ ) );
NOR3_X1 \malu/Shift/_1079_ ( .A1(\malu/Shift/_0135_ ), .A2(\malu/Shift/_0718_ ), .A3(\malu/Shift/_0717_ ), .ZN(\malu/Shift/_0325_ ) );
NOR3_X1 \malu/Shift/_1080_ ( .A1(\malu/Shift/_0325_ ), .A2(\malu/Shift/_0137_ ), .A3(\malu/Shift/_0253_ ), .ZN(\malu/Shift/_0326_ ) );
MUX2_X2 \malu/Shift/_1081_ ( .A(\malu/Shift/_0326_ ), .B(\malu/Shift/_0322_ ), .S(\malu/Shift/_0710_ ), .Z(\malu/Shift/_0327_ ) );
OAI21_X2 \malu/Shift/_1082_ ( .A(\malu/Shift/_0324_ ), .B1(\malu/Shift/_0327_ ), .B2(\malu/Shift/_0308_ ), .ZN(\malu/Shift/_0328_ ) );
NAND2_X1 \malu/Shift/_1083_ ( .A1(\malu/Shift/_0328_ ), .A2(\malu/Shift/_0720_ ), .ZN(\malu/Shift/_0329_ ) );
AND3_X1 \malu/Shift/_1084_ ( .A1(\malu/Shift/_0163_ ), .A2(\malu/Shift/_0168_ ), .A3(\malu/Shift/_0151_ ), .ZN(\malu/Shift/_0330_ ) );
AOI21_X1 \malu/Shift/_1085_ ( .A(\malu/Shift/_0100_ ), .B1(\malu/Shift/_0185_ ), .B2(\malu/Shift/_0189_ ), .ZN(\malu/Shift/_0331_ ) );
NOR3_X1 \malu/Shift/_1086_ ( .A1(\malu/Shift/_0330_ ), .A2(\malu/Shift/_0719_ ), .A3(\malu/Shift/_0331_ ), .ZN(\malu/Shift/_0332_ ) );
INV_X1 \malu/Shift/_1087_ ( .A(\malu/Shift/_0656_ ), .ZN(\malu/Shift/_0333_ ) );
NOR3_X1 \malu/Shift/_1088_ ( .A1(\malu/Shift/_0332_ ), .A2(\malu/Shift/_0720_ ), .A3(\malu/Shift/_0333_ ), .ZN(\malu/Shift/_0334_ ) );
BUF_X4 \malu/Shift/_1089_ ( .A(\malu/Shift/_0048_ ), .Z(\malu/Shift/_0335_ ) );
NAND3_X1 \malu/Shift/_1090_ ( .A1(\malu/Shift/_0118_ ), .A2(\malu/Shift/_0123_ ), .A3(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0336_ ) );
NAND3_X1 \malu/Shift/_1091_ ( .A1(\malu/Shift/_0174_ ), .A2(\malu/Shift/_0180_ ), .A3(\malu/Shift/_0151_ ), .ZN(\malu/Shift/_0337_ ) );
NAND2_X1 \malu/Shift/_1092_ ( .A1(\malu/Shift/_0336_ ), .A2(\malu/Shift/_0337_ ), .ZN(\malu/Shift/_0338_ ) );
OAI21_X1 \malu/Shift/_1093_ ( .A(\malu/Shift/_0334_ ), .B1(\malu/Shift/_0335_ ), .B2(\malu/Shift/_0338_ ), .ZN(\malu/Shift/_0339_ ) );
NAND3_X1 \malu/Shift/_1094_ ( .A1(\malu/Shift/_0714_ ), .A2(\malu/Shift/_0715_ ), .A3(\malu/Shift/_0027_ ), .ZN(\malu/Shift/_0340_ ) );
NOR2_X1 \malu/Shift/_1095_ ( .A1(\malu/Shift/_0202_ ), .A2(\malu/Shift/_0717_ ), .ZN(\malu/Shift/_0341_ ) );
OAI21_X1 \malu/Shift/_1096_ ( .A(\malu/Shift/_0033_ ), .B1(\malu/Shift/_0164_ ), .B2(\malu/Shift/_0157_ ), .ZN(\malu/Shift/_0342_ ) );
OAI21_X1 \malu/Shift/_1097_ ( .A(\malu/Shift/_0717_ ), .B1(\malu/Shift/_0156_ ), .B2(\malu/Shift/_0154_ ), .ZN(\malu/Shift/_0343_ ) );
NAND2_X1 \malu/Shift/_1098_ ( .A1(\malu/Shift/_0342_ ), .A2(\malu/Shift/_0343_ ), .ZN(\malu/Shift/_0344_ ) );
MUX2_X1 \malu/Shift/_1099_ ( .A(\malu/Shift/_0341_ ), .B(\malu/Shift/_0344_ ), .S(\malu/Shift/_0080_ ), .Z(\malu/Shift/_0345_ ) );
NAND3_X1 \malu/Shift/_1100_ ( .A1(\malu/Shift/_0345_ ), .A2(\malu/Shift/_0335_ ), .A3(\malu/Shift/_0205_ ), .ZN(\malu/Shift/_0346_ ) );
NAND4_X1 \malu/Shift/_1101_ ( .A1(\malu/Shift/_0329_ ), .A2(\malu/Shift/_0339_ ), .A3(\malu/Shift/_0340_ ), .A4(\malu/Shift/_0346_ ), .ZN(\malu/Shift/_0748_ ) );
MUX2_X1 \malu/Shift/_1102_ ( .A(\malu/Shift/_0219_ ), .B(\malu/Shift/_0214_ ), .S(\malu/Shift/_0051_ ), .Z(\malu/Shift/_0347_ ) );
NOR2_X1 \malu/Shift/_1103_ ( .A1(\malu/Shift/_0347_ ), .A2(\malu/Shift/_0719_ ), .ZN(\malu/Shift/_0348_ ) );
NOR4_X1 \malu/Shift/_1104_ ( .A1(\malu/Shift/_0098_ ), .A2(\malu/Shift/_0718_ ), .A3(\malu/Shift/_0717_ ), .A4(\malu/Shift/_0047_ ), .ZN(\malu/Shift/_0349_ ) );
OAI21_X1 \malu/Shift/_1105_ ( .A(\malu/Shift/_0194_ ), .B1(\malu/Shift/_0348_ ), .B2(\malu/Shift/_0349_ ), .ZN(\malu/Shift/_0350_ ) );
NOR2_X1 \malu/Shift/_1106_ ( .A1(\malu/Shift/_0098_ ), .A2(\malu/Shift/_0717_ ), .ZN(\malu/Shift/_0351_ ) );
AND2_X1 \malu/Shift/_1107_ ( .A1(\malu/Shift/_0351_ ), .A2(\malu/Shift/_0049_ ), .ZN(\malu/Shift/_0352_ ) );
NOR3_X1 \malu/Shift/_1108_ ( .A1(\malu/Shift/_0352_ ), .A2(\malu/Shift/_0137_ ), .A3(\malu/Shift/_0253_ ), .ZN(\malu/Shift/_0353_ ) );
MUX2_X2 \malu/Shift/_1109_ ( .A(\malu/Shift/_0353_ ), .B(\malu/Shift/_0347_ ), .S(\malu/Shift/_0711_ ), .Z(\malu/Shift/_0354_ ) );
OAI21_X1 \malu/Shift/_1110_ ( .A(\malu/Shift/_0350_ ), .B1(\malu/Shift/_0354_ ), .B2(\malu/Shift/_0308_ ), .ZN(\malu/Shift/_0355_ ) );
NAND2_X1 \malu/Shift/_1111_ ( .A1(\malu/Shift/_0355_ ), .A2(\malu/Shift/_0720_ ), .ZN(\malu/Shift/_0356_ ) );
AND3_X1 \malu/Shift/_1112_ ( .A1(\malu/Shift/_0207_ ), .A2(\malu/Shift/_0209_ ), .A3(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0357_ ) );
AOI21_X1 \malu/Shift/_1113_ ( .A(\malu/Shift/_0718_ ), .B1(\malu/Shift/_0229_ ), .B2(\malu/Shift/_0230_ ), .ZN(\malu/Shift/_0358_ ) );
OR2_X1 \malu/Shift/_1114_ ( .A1(\malu/Shift/_0357_ ), .A2(\malu/Shift/_0358_ ), .ZN(\malu/Shift/_0359_ ) );
AND2_X1 \malu/Shift/_1115_ ( .A1(\malu/Shift/_0226_ ), .A2(\malu/Shift/_0227_ ), .ZN(\malu/Shift/_0360_ ) );
MUX2_X2 \malu/Shift/_1116_ ( .A(\malu/Shift/_0239_ ), .B(\malu/Shift/_0360_ ), .S(\malu/Shift/_0718_ ), .Z(\malu/Shift/_0361_ ) );
MUX2_X2 \malu/Shift/_1117_ ( .A(\malu/Shift/_0359_ ), .B(\malu/Shift/_0361_ ), .S(\malu/Shift/_0064_ ), .Z(\malu/Shift/_0362_ ) );
AND2_X1 \malu/Shift/_1118_ ( .A1(\malu/Shift/_0656_ ), .A2(\malu/Shift/_0108_ ), .ZN(\malu/Shift/_0363_ ) );
OR3_X2 \malu/Shift/_1119_ ( .A1(\malu/Shift/_0054_ ), .A2(\malu/Shift/_0044_ ), .A3(\malu/Shift/_0693_ ), .ZN(\malu/Shift/_0364_ ) );
OR3_X1 \malu/Shift/_1120_ ( .A1(\malu/Shift/_0058_ ), .A2(\malu/Shift/_0055_ ), .A3(\malu/Shift/_0717_ ), .ZN(\malu/Shift/_0365_ ) );
NAND3_X1 \malu/Shift/_1121_ ( .A1(\malu/Shift/_0364_ ), .A2(\malu/Shift/_0365_ ), .A3(\malu/Shift/_0051_ ), .ZN(\malu/Shift/_0366_ ) );
OAI21_X1 \malu/Shift/_1122_ ( .A(\malu/Shift/_0366_ ), .B1(\malu/Shift/_0247_ ), .B2(\malu/Shift/_0080_ ), .ZN(\malu/Shift/_0367_ ) );
AND2_X1 \malu/Shift/_1123_ ( .A1(\malu/Shift/_0367_ ), .A2(\malu/Shift/_0047_ ), .ZN(\malu/Shift/_0368_ ) );
AOI22_X2 \malu/Shift/_1124_ ( .A1(\malu/Shift/_0362_ ), .A2(\malu/Shift/_0363_ ), .B1(\malu/Shift/_0205_ ), .B2(\malu/Shift/_0368_ ), .ZN(\malu/Shift/_0369_ ) );
OAI211_X2 \malu/Shift/_1125_ ( .A(\malu/Shift/_0356_ ), .B(\malu/Shift/_0369_ ), .C1(\malu/Shift/_0057_ ), .C2(\malu/Shift/_0105_ ), .ZN(\malu/Shift/_0749_ ) );
AOI21_X1 \malu/Shift/_1126_ ( .A(\malu/Shift/_0718_ ), .B1(\malu/Shift/_0256_ ), .B2(\malu/Shift/_0257_ ), .ZN(\malu/Shift/_0370_ ) );
AOI21_X1 \malu/Shift/_1127_ ( .A(\malu/Shift/_0370_ ), .B1(\malu/Shift/_0718_ ), .B2(\malu/Shift/_0251_ ), .ZN(\malu/Shift/_0371_ ) );
AND2_X1 \malu/Shift/_1128_ ( .A1(\malu/Shift/_0371_ ), .A2(\malu/Shift/_0711_ ), .ZN(\malu/Shift/_0372_ ) );
AND4_X1 \malu/Shift/_1129_ ( .A1(\malu/Shift/_0151_ ), .A2(\malu/Shift/_0197_ ), .A3(\malu/Shift/_0039_ ), .A4(\malu/Shift/_0719_ ), .ZN(\malu/Shift/_0373_ ) );
OAI21_X1 \malu/Shift/_1130_ ( .A(\malu/Shift/_0194_ ), .B1(\malu/Shift/_0372_ ), .B2(\malu/Shift/_0373_ ), .ZN(\malu/Shift/_0374_ ) );
AND2_X1 \malu/Shift/_1131_ ( .A1(\malu/Shift/_0719_ ), .A2(\malu/Shift/_0024_ ), .ZN(\malu/Shift/_0375_ ) );
OAI21_X1 \malu/Shift/_1132_ ( .A(\malu/Shift/_0113_ ), .B1(\malu/Shift/_0372_ ), .B2(\malu/Shift/_0375_ ), .ZN(\malu/Shift/_0376_ ) );
NAND2_X1 \malu/Shift/_1133_ ( .A1(\malu/Shift/_0374_ ), .A2(\malu/Shift/_0376_ ), .ZN(\malu/Shift/_0377_ ) );
NAND2_X1 \malu/Shift/_1134_ ( .A1(\malu/Shift/_0377_ ), .A2(\malu/Shift/_0720_ ), .ZN(\malu/Shift/_0378_ ) );
NAND2_X1 \malu/Shift/_1135_ ( .A1(\malu/Shift/_0273_ ), .A2(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0379_ ) );
OAI211_X2 \malu/Shift/_1136_ ( .A(\malu/Shift/_0379_ ), .B(\malu/Shift/_0048_ ), .C1(\malu/Shift/_0269_ ), .C2(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0380_ ) );
NAND3_X1 \malu/Shift/_1137_ ( .A1(\malu/Shift/_0259_ ), .A2(\malu/Shift/_0260_ ), .A3(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0381_ ) );
NAND3_X1 \malu/Shift/_1138_ ( .A1(\malu/Shift/_0275_ ), .A2(\malu/Shift/_0053_ ), .A3(\malu/Shift/_0276_ ), .ZN(\malu/Shift/_0382_ ) );
NAND3_X1 \malu/Shift/_1139_ ( .A1(\malu/Shift/_0381_ ), .A2(\malu/Shift/_0382_ ), .A3(\malu/Shift/_0719_ ), .ZN(\malu/Shift/_0383_ ) );
NAND3_X1 \malu/Shift/_1140_ ( .A1(\malu/Shift/_0380_ ), .A2(\malu/Shift/_0363_ ), .A3(\malu/Shift/_0383_ ), .ZN(\malu/Shift/_0384_ ) );
NAND3_X1 \malu/Shift/_1141_ ( .A1(\malu/Shift/_0714_ ), .A2(\malu/Shift/_0715_ ), .A3(\malu/Shift/_0029_ ), .ZN(\malu/Shift/_0385_ ) );
OAI21_X1 \malu/Shift/_1142_ ( .A(\malu/Shift/_0033_ ), .B1(\malu/Shift/_0161_ ), .B2(\malu/Shift/_0166_ ), .ZN(\malu/Shift/_0386_ ) );
OAI21_X1 \malu/Shift/_1143_ ( .A(\malu/Shift/_0717_ ), .B1(\malu/Shift/_0164_ ), .B2(\malu/Shift/_0157_ ), .ZN(\malu/Shift/_0387_ ) );
NAND2_X1 \malu/Shift/_1144_ ( .A1(\malu/Shift/_0386_ ), .A2(\malu/Shift/_0387_ ), .ZN(\malu/Shift/_0388_ ) );
NAND2_X1 \malu/Shift/_1145_ ( .A1(\malu/Shift/_0388_ ), .A2(\malu/Shift/_0053_ ), .ZN(\malu/Shift/_0389_ ) );
OAI21_X1 \malu/Shift/_1146_ ( .A(\malu/Shift/_0389_ ), .B1(\malu/Shift/_0288_ ), .B2(\malu/Shift/_0053_ ), .ZN(\malu/Shift/_0390_ ) );
NAND3_X1 \malu/Shift/_1147_ ( .A1(\malu/Shift/_0390_ ), .A2(\malu/Shift/_0335_ ), .A3(\malu/Shift/_0205_ ), .ZN(\malu/Shift/_0391_ ) );
NAND4_X1 \malu/Shift/_1148_ ( .A1(\malu/Shift/_0378_ ), .A2(\malu/Shift/_0384_ ), .A3(\malu/Shift/_0385_ ), .A4(\malu/Shift/_0391_ ), .ZN(\malu/Shift/_0750_ ) );
OR2_X1 \malu/Shift/_1149_ ( .A1(\malu/Shift/_0099_ ), .A2(\malu/Shift/_0051_ ), .ZN(\malu/Shift/_0392_ ) );
NAND2_X1 \malu/Shift/_1150_ ( .A1(\malu/Shift/_0392_ ), .A2(\malu/Shift/_0091_ ), .ZN(\malu/Shift/_0393_ ) );
AND2_X1 \malu/Shift/_1151_ ( .A1(\malu/Shift/_0393_ ), .A2(\malu/Shift/_0711_ ), .ZN(\malu/Shift/_0394_ ) );
OAI21_X1 \malu/Shift/_1152_ ( .A(\malu/Shift/_0113_ ), .B1(\malu/Shift/_0394_ ), .B2(\malu/Shift/_0375_ ), .ZN(\malu/Shift/_0395_ ) );
AND2_X2 \malu/Shift/_1153_ ( .A1(\malu/Shift/_0194_ ), .A2(\malu/Shift/_0710_ ), .ZN(\malu/Shift/_0396_ ) );
NAND2_X1 \malu/Shift/_1154_ ( .A1(\malu/Shift/_0393_ ), .A2(\malu/Shift/_0396_ ), .ZN(\malu/Shift/_0397_ ) );
AND3_X1 \malu/Shift/_1155_ ( .A1(\malu/Shift/_0395_ ), .A2(\malu/Shift/_0720_ ), .A3(\malu/Shift/_0397_ ), .ZN(\malu/Shift/_0398_ ) );
OAI21_X1 \malu/Shift/_1156_ ( .A(\malu/Shift/_0719_ ), .B1(\malu/Shift/_0072_ ), .B2(\malu/Shift/_0081_ ), .ZN(\malu/Shift/_0399_ ) );
OAI21_X1 \malu/Shift/_1157_ ( .A(\malu/Shift/_0236_ ), .B1(\malu/Shift/_0699_ ), .B2(\malu/Shift/_0709_ ), .ZN(\malu/Shift/_0400_ ) );
NAND3_X1 \malu/Shift/_1158_ ( .A1(\malu/Shift/_0399_ ), .A2(\malu/Shift/_0400_ ), .A3(\malu/Shift/_0656_ ), .ZN(\malu/Shift/_0401_ ) );
INV_X1 \malu/Shift/_1159_ ( .A(\malu/Shift/_0646_ ), .ZN(\malu/Shift/_0402_ ) );
INV_X1 \malu/Shift/_1160_ ( .A(\malu/Shift/_0106_ ), .ZN(\malu/Shift/_0403_ ) );
AOI21_X1 \malu/Shift/_1161_ ( .A(\malu/Shift/_0402_ ), .B1(\malu/Shift/_0403_ ), .B2(\malu/Shift/_0719_ ), .ZN(\malu/Shift/_0404_ ) );
NAND2_X1 \malu/Shift/_1162_ ( .A1(\malu/Shift/_0295_ ), .A2(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0405_ ) );
OR3_X1 \malu/Shift/_1163_ ( .A1(\malu/Shift/_0058_ ), .A2(\malu/Shift/_0055_ ), .A3(\malu/Shift/_0693_ ), .ZN(\malu/Shift/_0406_ ) );
OR3_X1 \malu/Shift/_1164_ ( .A1(\malu/Shift/_0696_ ), .A2(\malu/Shift/_0059_ ), .A3(\malu/Shift/_0717_ ), .ZN(\malu/Shift/_0407_ ) );
NAND3_X1 \malu/Shift/_1165_ ( .A1(\malu/Shift/_0406_ ), .A2(\malu/Shift/_0407_ ), .A3(\malu/Shift/_0151_ ), .ZN(\malu/Shift/_0408_ ) );
NAND2_X1 \malu/Shift/_1166_ ( .A1(\malu/Shift/_0405_ ), .A2(\malu/Shift/_0408_ ), .ZN(\malu/Shift/_0409_ ) );
OAI21_X1 \malu/Shift/_1167_ ( .A(\malu/Shift/_0404_ ), .B1(\malu/Shift/_0409_ ), .B2(\malu/Shift/_0719_ ), .ZN(\malu/Shift/_0410_ ) );
AND3_X1 \malu/Shift/_1168_ ( .A1(\malu/Shift/_0401_ ), .A2(\malu/Shift/_0148_ ), .A3(\malu/Shift/_0410_ ), .ZN(\malu/Shift/_0411_ ) );
OAI22_X1 \malu/Shift/_1169_ ( .A1(\malu/Shift/_0398_ ), .A2(\malu/Shift/_0411_ ), .B1(\malu/Shift/_0695_ ), .B2(\malu/Shift/_0105_ ), .ZN(\malu/Shift/_0751_ ) );
AOI21_X1 \malu/Shift/_1170_ ( .A(\malu/Shift/_0333_ ), .B1(\malu/Shift/_0132_ ), .B2(\malu/Shift/_0719_ ), .ZN(\malu/Shift/_0412_ ) );
OAI21_X1 \malu/Shift/_1171_ ( .A(\malu/Shift/_0047_ ), .B1(\malu/Shift/_0181_ ), .B2(\malu/Shift/_0190_ ), .ZN(\malu/Shift/_0413_ ) );
NAND3_X1 \malu/Shift/_1172_ ( .A1(\malu/Shift/_0342_ ), .A2(\malu/Shift/_0343_ ), .A3(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0414_ ) );
OR3_X4 \malu/Shift/_1173_ ( .A1(\malu/Shift/_0161_ ), .A2(\malu/Shift/_0692_ ), .A3(\malu/Shift/_0166_ ), .ZN(\malu/Shift/_0415_ ) );
INV_X1 \malu/Shift/_1174_ ( .A(\malu/Shift/_0162_ ), .ZN(\malu/Shift/_0416_ ) );
OAI211_X2 \malu/Shift/_1175_ ( .A(\malu/Shift/_0416_ ), .B(\malu/Shift/_0692_ ), .C1(\malu/Shift/_0716_ ), .C2(\malu/Shift/_0182_ ), .ZN(\malu/Shift/_0417_ ) );
AND2_X4 \malu/Shift/_1176_ ( .A1(\malu/Shift/_0415_ ), .A2(\malu/Shift/_0417_ ), .ZN(\malu/Shift/_0418_ ) );
OR2_X4 \malu/Shift/_1177_ ( .A1(\malu/Shift/_0418_ ), .A2(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0419_ ) );
AND2_X4 \malu/Shift/_1178_ ( .A1(\malu/Shift/_0414_ ), .A2(\malu/Shift/_0419_ ), .ZN(\malu/Shift/_0420_ ) );
MUX2_X2 \malu/Shift/_1179_ ( .A(\malu/Shift/_0203_ ), .B(\malu/Shift/_0420_ ), .S(\malu/Shift/_0710_ ), .Z(\malu/Shift/_0421_ ) );
AOI221_X2 \malu/Shift/_1180_ ( .A(\malu/Shift/_0720_ ), .B1(\malu/Shift/_0412_ ), .B2(\malu/Shift/_0413_ ), .C1(\malu/Shift/_0249_ ), .C2(\malu/Shift/_0421_ ), .ZN(\malu/Shift/_0422_ ) );
NAND2_X1 \malu/Shift/_1181_ ( .A1(\malu/Shift/_0146_ ), .A2(\malu/Shift/_0048_ ), .ZN(\malu/Shift/_0423_ ) );
INV_X1 \malu/Shift/_1182_ ( .A(\malu/Shift/_0375_ ), .ZN(\malu/Shift/_0424_ ) );
AOI21_X1 \malu/Shift/_1183_ ( .A(\malu/Shift/_0308_ ), .B1(\malu/Shift/_0423_ ), .B2(\malu/Shift/_0424_ ), .ZN(\malu/Shift/_0425_ ) );
INV_X1 \malu/Shift/_1184_ ( .A(\malu/Shift/_0396_ ), .ZN(\malu/Shift/_0426_ ) );
NOR2_X1 \malu/Shift/_1185_ ( .A1(\malu/Shift/_0199_ ), .A2(\malu/Shift/_0426_ ), .ZN(\malu/Shift/_0427_ ) );
NOR3_X1 \malu/Shift/_1186_ ( .A1(\malu/Shift/_0425_ ), .A2(\malu/Shift/_0149_ ), .A3(\malu/Shift/_0427_ ), .ZN(\malu/Shift/_0428_ ) );
OAI22_X1 \malu/Shift/_1187_ ( .A1(\malu/Shift/_0422_ ), .A2(\malu/Shift/_0428_ ), .B1(\malu/Shift/_0182_ ), .B2(\malu/Shift/_0105_ ), .ZN(\malu/Shift/_0752_ ) );
AOI21_X1 \malu/Shift/_1188_ ( .A(\malu/Shift/_0375_ ), .B1(\malu/Shift/_0223_ ), .B2(\malu/Shift/_0711_ ), .ZN(\malu/Shift/_0429_ ) );
OR2_X1 \malu/Shift/_1189_ ( .A1(\malu/Shift/_0429_ ), .A2(\malu/Shift/_0308_ ), .ZN(\malu/Shift/_0430_ ) );
AND2_X1 \malu/Shift/_1190_ ( .A1(\malu/Shift/_0220_ ), .A2(\malu/Shift/_0222_ ), .ZN(\malu/Shift/_0431_ ) );
OR2_X1 \malu/Shift/_1191_ ( .A1(\malu/Shift/_0431_ ), .A2(\malu/Shift/_0426_ ), .ZN(\malu/Shift/_0432_ ) );
AND3_X1 \malu/Shift/_1192_ ( .A1(\malu/Shift/_0430_ ), .A2(\malu/Shift/_0720_ ), .A3(\malu/Shift/_0432_ ), .ZN(\malu/Shift/_0433_ ) );
NOR3_X1 \malu/Shift/_1193_ ( .A1(\malu/Shift/_0247_ ), .A2(\malu/Shift/_0718_ ), .A3(\malu/Shift/_0710_ ), .ZN(\malu/Shift/_0434_ ) );
NAND3_X1 \malu/Shift/_1194_ ( .A1(\malu/Shift/_0364_ ), .A2(\malu/Shift/_0365_ ), .A3(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0435_ ) );
OR3_X1 \malu/Shift/_1195_ ( .A1(\malu/Shift/_0696_ ), .A2(\malu/Shift/_0059_ ), .A3(\malu/Shift/_0693_ ), .ZN(\malu/Shift/_0436_ ) );
OR3_X1 \malu/Shift/_1196_ ( .A1(\malu/Shift/_0676_ ), .A2(\malu/Shift/_0697_ ), .A3(\malu/Shift/_0717_ ), .ZN(\malu/Shift/_0437_ ) );
NAND3_X1 \malu/Shift/_1197_ ( .A1(\malu/Shift/_0436_ ), .A2(\malu/Shift/_0437_ ), .A3(\malu/Shift/_0050_ ), .ZN(\malu/Shift/_0438_ ) );
AOI21_X1 \malu/Shift/_1198_ ( .A(\malu/Shift/_0719_ ), .B1(\malu/Shift/_0435_ ), .B2(\malu/Shift/_0438_ ), .ZN(\malu/Shift/_0439_ ) );
OR2_X2 \malu/Shift/_1199_ ( .A1(\malu/Shift/_0434_ ), .A2(\malu/Shift/_0439_ ), .ZN(\malu/Shift/_0440_ ) );
MUX2_X1 \malu/Shift/_1200_ ( .A(\malu/Shift/_0232_ ), .B(\malu/Shift/_0215_ ), .S(\malu/Shift/_0719_ ), .Z(\malu/Shift/_0441_ ) );
AOI221_X2 \malu/Shift/_1201_ ( .A(\malu/Shift/_0720_ ), .B1(\malu/Shift/_0249_ ), .B2(\malu/Shift/_0440_ ), .C1(\malu/Shift/_0441_ ), .C2(\malu/Shift/_0656_ ), .ZN(\malu/Shift/_0442_ ) );
OAI22_X1 \malu/Shift/_1202_ ( .A1(\malu/Shift/_0433_ ), .A2(\malu/Shift/_0442_ ), .B1(\malu/Shift/_0666_ ), .B2(\malu/Shift/_0105_ ), .ZN(\malu/Shift/_0722_ ) );
AOI21_X1 \malu/Shift/_1203_ ( .A(\malu/Shift/_0719_ ), .B1(\malu/Shift/_0252_ ), .B2(\malu/Shift/_0254_ ), .ZN(\malu/Shift/_0443_ ) );
OAI21_X1 \malu/Shift/_1204_ ( .A(\malu/Shift/_0112_ ), .B1(\malu/Shift/_0443_ ), .B2(\malu/Shift/_0375_ ), .ZN(\malu/Shift/_0444_ ) );
NAND2_X1 \malu/Shift/_1205_ ( .A1(\malu/Shift/_0284_ ), .A2(\malu/Shift/_0396_ ), .ZN(\malu/Shift/_0445_ ) );
AND3_X1 \malu/Shift/_1206_ ( .A1(\malu/Shift/_0444_ ), .A2(\malu/Shift/_0720_ ), .A3(\malu/Shift/_0445_ ), .ZN(\malu/Shift/_0446_ ) );
NAND3_X1 \malu/Shift/_1207_ ( .A1(\malu/Shift/_0258_ ), .A2(\malu/Shift/_0261_ ), .A3(\malu/Shift/_0719_ ), .ZN(\malu/Shift/_0447_ ) );
AND2_X1 \malu/Shift/_1208_ ( .A1(\malu/Shift/_0447_ ), .A2(\malu/Shift/_0656_ ), .ZN(\malu/Shift/_0448_ ) );
NAND3_X1 \malu/Shift/_1209_ ( .A1(\malu/Shift/_0274_ ), .A2(\malu/Shift/_0277_ ), .A3(\malu/Shift/_0047_ ), .ZN(\malu/Shift/_0449_ ) );
OR3_X1 \malu/Shift/_1210_ ( .A1(\malu/Shift/_0288_ ), .A2(\malu/Shift/_0718_ ), .A3(\malu/Shift/_0710_ ), .ZN(\malu/Shift/_0450_ ) );
NAND2_X1 \malu/Shift/_1211_ ( .A1(\malu/Shift/_0388_ ), .A2(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0451_ ) );
OR3_X4 \malu/Shift/_1212_ ( .A1(\malu/Shift/_0187_ ), .A2(\malu/Shift/_0184_ ), .A3(\malu/Shift/_0717_ ), .ZN(\malu/Shift/_0452_ ) );
OAI211_X2 \malu/Shift/_1213_ ( .A(\malu/Shift/_0416_ ), .B(\malu/Shift/_0717_ ), .C1(\malu/Shift/_0716_ ), .C2(\malu/Shift/_0182_ ), .ZN(\malu/Shift/_0453_ ) );
NAND3_X1 \malu/Shift/_1214_ ( .A1(\malu/Shift/_0452_ ), .A2(\malu/Shift/_0453_ ), .A3(\malu/Shift/_0051_ ), .ZN(\malu/Shift/_0454_ ) );
NAND2_X1 \malu/Shift/_1215_ ( .A1(\malu/Shift/_0451_ ), .A2(\malu/Shift/_0454_ ), .ZN(\malu/Shift/_0455_ ) );
NAND2_X1 \malu/Shift/_1216_ ( .A1(\malu/Shift/_0455_ ), .A2(\malu/Shift/_0047_ ), .ZN(\malu/Shift/_0456_ ) );
NAND2_X1 \malu/Shift/_1217_ ( .A1(\malu/Shift/_0450_ ), .A2(\malu/Shift/_0456_ ), .ZN(\malu/Shift/_0457_ ) );
AOI221_X1 \malu/Shift/_1218_ ( .A(\malu/Shift/_0720_ ), .B1(\malu/Shift/_0448_ ), .B2(\malu/Shift/_0449_ ), .C1(\malu/Shift/_0249_ ), .C2(\malu/Shift/_0457_ ), .ZN(\malu/Shift/_0458_ ) );
OAI22_X1 \malu/Shift/_1219_ ( .A1(\malu/Shift/_0446_ ), .A2(\malu/Shift/_0458_ ), .B1(\malu/Shift/_0186_ ), .B2(\malu/Shift/_0105_ ), .ZN(\malu/Shift/_0723_ ) );
OR3_X1 \malu/Shift/_1220_ ( .A1(\malu/Shift/_0676_ ), .A2(\malu/Shift/_0697_ ), .A3(\malu/Shift/_0693_ ), .ZN(\malu/Shift/_0459_ ) );
OR3_X1 \malu/Shift/_1221_ ( .A1(\malu/Shift/_0702_ ), .A2(\malu/Shift/_0686_ ), .A3(\malu/Shift/_0717_ ), .ZN(\malu/Shift/_0460_ ) );
NAND3_X1 \malu/Shift/_1222_ ( .A1(\malu/Shift/_0459_ ), .A2(\malu/Shift/_0460_ ), .A3(\malu/Shift/_0050_ ), .ZN(\malu/Shift/_0461_ ) );
NAND3_X1 \malu/Shift/_1223_ ( .A1(\malu/Shift/_0406_ ), .A2(\malu/Shift/_0407_ ), .A3(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0462_ ) );
NAND2_X1 \malu/Shift/_1224_ ( .A1(\malu/Shift/_0461_ ), .A2(\malu/Shift/_0462_ ), .ZN(\malu/Shift/_0463_ ) );
MUX2_X1 \malu/Shift/_1225_ ( .A(\malu/Shift/_0463_ ), .B(\malu/Shift/_0298_ ), .S(\malu/Shift/_0719_ ), .Z(\malu/Shift/_0464_ ) );
MUX2_X1 \malu/Shift/_1226_ ( .A(\malu/Shift/_0302_ ), .B(\malu/Shift/_0313_ ), .S(\malu/Shift/_0719_ ), .Z(\malu/Shift/_0465_ ) );
AOI221_X1 \malu/Shift/_1227_ ( .A(\malu/Shift/_0720_ ), .B1(\malu/Shift/_0464_ ), .B2(\malu/Shift/_0646_ ), .C1(\malu/Shift/_0656_ ), .C2(\malu/Shift/_0465_ ), .ZN(\malu/Shift/_0466_ ) );
OAI21_X1 \malu/Shift/_1228_ ( .A(\malu/Shift/_0047_ ), .B1(\malu/Shift/_0309_ ), .B2(\malu/Shift/_0253_ ), .ZN(\malu/Shift/_0467_ ) );
NAND2_X1 \malu/Shift/_1229_ ( .A1(\malu/Shift/_0467_ ), .A2(\malu/Shift/_0424_ ), .ZN(\malu/Shift/_0468_ ) );
AOI221_X4 \malu/Shift/_1230_ ( .A(\malu/Shift/_0108_ ), .B1(\malu/Shift/_0309_ ), .B2(\malu/Shift/_0396_ ), .C1(\malu/Shift/_0468_ ), .C2(\malu/Shift/_0113_ ), .ZN(\malu/Shift/_0469_ ) );
OAI22_X1 \malu/Shift/_1231_ ( .A1(\malu/Shift/_0466_ ), .A2(\malu/Shift/_0469_ ), .B1(\malu/Shift/_0701_ ), .B2(\malu/Shift/_0105_ ), .ZN(\malu/Shift/_0724_ ) );
AOI21_X1 \malu/Shift/_1232_ ( .A(\malu/Shift/_0333_ ), .B1(\malu/Shift/_0322_ ), .B2(\malu/Shift/_0719_ ), .ZN(\malu/Shift/_0470_ ) );
OAI21_X1 \malu/Shift/_1233_ ( .A(\malu/Shift/_0470_ ), .B1(\malu/Shift/_0719_ ), .B2(\malu/Shift/_0338_ ), .ZN(\malu/Shift/_0471_ ) );
NAND2_X1 \malu/Shift/_1234_ ( .A1(\malu/Shift/_0345_ ), .A2(\malu/Shift/_0719_ ), .ZN(\malu/Shift/_0472_ ) );
OAI21_X1 \malu/Shift/_1235_ ( .A(\malu/Shift/_0034_ ), .B1(\malu/Shift/_0172_ ), .B2(\malu/Shift/_0188_ ), .ZN(\malu/Shift/_0473_ ) );
OAI21_X1 \malu/Shift/_1236_ ( .A(\malu/Shift/_0717_ ), .B1(\malu/Shift/_0187_ ), .B2(\malu/Shift/_0184_ ), .ZN(\malu/Shift/_0474_ ) );
NAND3_X1 \malu/Shift/_1237_ ( .A1(\malu/Shift/_0473_ ), .A2(\malu/Shift/_0474_ ), .A3(\malu/Shift/_0080_ ), .ZN(\malu/Shift/_0475_ ) );
OAI211_X2 \malu/Shift/_1238_ ( .A(\malu/Shift/_0711_ ), .B(\malu/Shift/_0475_ ), .C1(\malu/Shift/_0418_ ), .C2(\malu/Shift/_0100_ ), .ZN(\malu/Shift/_0476_ ) );
NAND2_X1 \malu/Shift/_1239_ ( .A1(\malu/Shift/_0472_ ), .A2(\malu/Shift/_0476_ ), .ZN(\malu/Shift/_0477_ ) );
NAND2_X1 \malu/Shift/_1240_ ( .A1(\malu/Shift/_0477_ ), .A2(\malu/Shift/_0249_ ), .ZN(\malu/Shift/_0478_ ) );
NAND3_X1 \malu/Shift/_1241_ ( .A1(\malu/Shift/_0471_ ), .A2(\malu/Shift/_0148_ ), .A3(\malu/Shift/_0478_ ), .ZN(\malu/Shift/_0479_ ) );
OR3_X1 \malu/Shift/_1242_ ( .A1(\malu/Shift/_0198_ ), .A2(\malu/Shift/_0718_ ), .A3(\malu/Shift/_0426_ ), .ZN(\malu/Shift/_0480_ ) );
MUX2_X1 \malu/Shift/_1243_ ( .A(\malu/Shift/_0097_ ), .B(\malu/Shift/_0326_ ), .S(\malu/Shift/_0711_ ), .Z(\malu/Shift/_0481_ ) );
OAI21_X1 \malu/Shift/_1244_ ( .A(\malu/Shift/_0480_ ), .B1(\malu/Shift/_0481_ ), .B2(\malu/Shift/_0308_ ), .ZN(\malu/Shift/_0482_ ) );
OAI21_X1 \malu/Shift/_1245_ ( .A(\malu/Shift/_0479_ ), .B1(\malu/Shift/_0149_ ), .B2(\malu/Shift/_0482_ ), .ZN(\malu/Shift/_0483_ ) );
OAI21_X1 \malu/Shift/_1246_ ( .A(\malu/Shift/_0483_ ), .B1(\malu/Shift/_0171_ ), .B2(\malu/Shift/_0105_ ), .ZN(\malu/Shift/_0725_ ) );
AOI21_X1 \malu/Shift/_1247_ ( .A(\malu/Shift/_0333_ ), .B1(\malu/Shift/_0347_ ), .B2(\malu/Shift/_0719_ ), .ZN(\malu/Shift/_0484_ ) );
OR3_X4 \malu/Shift/_1248_ ( .A1(\malu/Shift/_0357_ ), .A2(\malu/Shift/_0719_ ), .A3(\malu/Shift/_0358_ ), .ZN(\malu/Shift/_0485_ ) );
AOI21_X2 \malu/Shift/_1249_ ( .A(\malu/Shift/_0051_ ), .B1(\malu/Shift/_0436_ ), .B2(\malu/Shift/_0437_ ), .ZN(\malu/Shift/_0486_ ) );
OR3_X2 \malu/Shift/_1250_ ( .A1(\malu/Shift/_0702_ ), .A2(\malu/Shift/_0686_ ), .A3(\malu/Shift/_0693_ ), .ZN(\malu/Shift/_0487_ ) );
OR3_X2 \malu/Shift/_1251_ ( .A1(\malu/Shift/_0706_ ), .A2(\malu/Shift/_0703_ ), .A3(\malu/Shift/_0717_ ), .ZN(\malu/Shift/_0488_ ) );
AOI21_X2 \malu/Shift/_1252_ ( .A(\malu/Shift/_0718_ ), .B1(\malu/Shift/_0487_ ), .B2(\malu/Shift/_0488_ ), .ZN(\malu/Shift/_0489_ ) );
NOR2_X2 \malu/Shift/_1253_ ( .A1(\malu/Shift/_0486_ ), .A2(\malu/Shift/_0489_ ), .ZN(\malu/Shift/_0490_ ) );
MUX2_X2 \malu/Shift/_1254_ ( .A(\malu/Shift/_0490_ ), .B(\malu/Shift/_0367_ ), .S(\malu/Shift/_0719_ ), .Z(\malu/Shift/_0491_ ) );
AOI221_X1 \malu/Shift/_1255_ ( .A(\malu/Shift/_0720_ ), .B1(\malu/Shift/_0484_ ), .B2(\malu/Shift/_0485_ ), .C1(\malu/Shift/_0249_ ), .C2(\malu/Shift/_0491_ ), .ZN(\malu/Shift/_0492_ ) );
OAI21_X1 \malu/Shift/_1256_ ( .A(\malu/Shift/_0424_ ), .B1(\malu/Shift/_0353_ ), .B2(\malu/Shift/_0719_ ), .ZN(\malu/Shift/_0493_ ) );
AOI221_X4 \malu/Shift/_1257_ ( .A(\malu/Shift/_0108_ ), .B1(\malu/Shift/_0352_ ), .B2(\malu/Shift/_0396_ ), .C1(\malu/Shift/_0493_ ), .C2(\malu/Shift/_0112_ ), .ZN(\malu/Shift/_0494_ ) );
OAI22_X1 \malu/Shift/_1258_ ( .A1(\malu/Shift/_0492_ ), .A2(\malu/Shift/_0494_ ), .B1(\malu/Shift/_0705_ ), .B2(\malu/Shift/_0105_ ), .ZN(\malu/Shift/_0726_ ) );
NAND3_X1 \malu/Shift/_1259_ ( .A1(\malu/Shift/_0381_ ), .A2(\malu/Shift/_0382_ ), .A3(\malu/Shift/_0048_ ), .ZN(\malu/Shift/_0495_ ) );
OAI211_X2 \malu/Shift/_1260_ ( .A(\malu/Shift/_0363_ ), .B(\malu/Shift/_0495_ ), .C1(\malu/Shift/_0371_ ), .C2(\malu/Shift/_0335_ ), .ZN(\malu/Shift/_0496_ ) );
OAI211_X2 \malu/Shift/_1261_ ( .A(\malu/Shift/_0389_ ), .B(\malu/Shift/_0719_ ), .C1(\malu/Shift/_0288_ ), .C2(\malu/Shift/_0053_ ), .ZN(\malu/Shift/_0497_ ) );
OAI21_X1 \malu/Shift/_1262_ ( .A(\malu/Shift/_0034_ ), .B1(\malu/Shift/_0176_ ), .B2(\malu/Shift/_0173_ ), .ZN(\malu/Shift/_0498_ ) );
OAI21_X1 \malu/Shift/_1263_ ( .A(\malu/Shift/_0717_ ), .B1(\malu/Shift/_0172_ ), .B2(\malu/Shift/_0188_ ), .ZN(\malu/Shift/_0499_ ) );
NAND2_X1 \malu/Shift/_1264_ ( .A1(\malu/Shift/_0498_ ), .A2(\malu/Shift/_0499_ ), .ZN(\malu/Shift/_0500_ ) );
NAND2_X1 \malu/Shift/_1265_ ( .A1(\malu/Shift/_0500_ ), .A2(\malu/Shift/_0100_ ), .ZN(\malu/Shift/_0501_ ) );
NAND3_X1 \malu/Shift/_1266_ ( .A1(\malu/Shift/_0452_ ), .A2(\malu/Shift/_0453_ ), .A3(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0502_ ) );
NAND3_X1 \malu/Shift/_1267_ ( .A1(\malu/Shift/_0501_ ), .A2(\malu/Shift/_0502_ ), .A3(\malu/Shift/_0048_ ), .ZN(\malu/Shift/_0503_ ) );
NAND3_X1 \malu/Shift/_1268_ ( .A1(\malu/Shift/_0497_ ), .A2(\malu/Shift/_0205_ ), .A3(\malu/Shift/_0503_ ), .ZN(\malu/Shift/_0504_ ) );
AND3_X1 \malu/Shift/_1269_ ( .A1(\malu/Shift/_0197_ ), .A2(\malu/Shift/_0053_ ), .A3(\malu/Shift/_0039_ ), .ZN(\malu/Shift/_0505_ ) );
NAND3_X1 \malu/Shift/_1270_ ( .A1(\malu/Shift/_0196_ ), .A2(\malu/Shift/_0505_ ), .A3(\malu/Shift/_0335_ ), .ZN(\malu/Shift/_0506_ ) );
AND2_X1 \malu/Shift/_1271_ ( .A1(\malu/Shift/_0720_ ), .A2(\malu/Shift/_0024_ ), .ZN(\malu/Shift/_0507_ ) );
AOI22_X1 \malu/Shift/_1272_ ( .A1(\malu/Shift/_0113_ ), .A2(\malu/Shift/_0507_ ), .B1(\malu/Shift/_0635_ ), .B2(\malu/Shift/_0006_ ), .ZN(\malu/Shift/_0508_ ) );
NAND4_X1 \malu/Shift/_1273_ ( .A1(\malu/Shift/_0496_ ), .A2(\malu/Shift/_0504_ ), .A3(\malu/Shift/_0506_ ), .A4(\malu/Shift/_0508_ ), .ZN(\malu/Shift/_0727_ ) );
AOI21_X1 \malu/Shift/_1274_ ( .A(\malu/Shift/_0402_ ), .B1(\malu/Shift/_0107_ ), .B2(\malu/Shift/_0720_ ), .ZN(\malu/Shift/_0509_ ) );
OR3_X1 \malu/Shift/_1275_ ( .A1(\malu/Shift/_0073_ ), .A2(\malu/Shift/_0707_ ), .A3(\malu/Shift/_0717_ ), .ZN(\malu/Shift/_0510_ ) );
OR3_X1 \malu/Shift/_1276_ ( .A1(\malu/Shift/_0706_ ), .A2(\malu/Shift/_0703_ ), .A3(\malu/Shift/_0038_ ), .ZN(\malu/Shift/_0511_ ) );
NAND3_X1 \malu/Shift/_1277_ ( .A1(\malu/Shift/_0510_ ), .A2(\malu/Shift/_0151_ ), .A3(\malu/Shift/_0511_ ), .ZN(\malu/Shift/_0512_ ) );
NAND3_X1 \malu/Shift/_1278_ ( .A1(\malu/Shift/_0459_ ), .A2(\malu/Shift/_0460_ ), .A3(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0513_ ) );
NAND2_X1 \malu/Shift/_1279_ ( .A1(\malu/Shift/_0512_ ), .A2(\malu/Shift/_0513_ ), .ZN(\malu/Shift/_0514_ ) );
MUX2_X1 \malu/Shift/_1280_ ( .A(\malu/Shift/_0514_ ), .B(\malu/Shift/_0409_ ), .S(\malu/Shift/_0719_ ), .Z(\malu/Shift/_0515_ ) );
OAI21_X1 \malu/Shift/_1281_ ( .A(\malu/Shift/_0509_ ), .B1(\malu/Shift/_0515_ ), .B2(\malu/Shift/_0720_ ), .ZN(\malu/Shift/_0516_ ) );
AND2_X1 \malu/Shift/_1282_ ( .A1(\malu/Shift/_0112_ ), .A2(\malu/Shift/_0507_ ), .ZN(\malu/Shift/_0517_ ) );
INV_X1 \malu/Shift/_1283_ ( .A(\malu/Shift/_0517_ ), .ZN(\malu/Shift/_0518_ ) );
NAND3_X1 \malu/Shift/_1284_ ( .A1(\malu/Shift/_0082_ ), .A2(\malu/Shift/_0101_ ), .A3(\malu/Shift/_0363_ ), .ZN(\malu/Shift/_0519_ ) );
NAND3_X1 \malu/Shift/_1285_ ( .A1(\malu/Shift/_0714_ ), .A2(\malu/Shift/_0715_ ), .A3(\malu/Shift/_0007_ ), .ZN(\malu/Shift/_0520_ ) );
NAND4_X1 \malu/Shift/_1286_ ( .A1(\malu/Shift/_0516_ ), .A2(\malu/Shift/_0518_ ), .A3(\malu/Shift/_0519_ ), .A4(\malu/Shift/_0520_ ), .ZN(\malu/Shift/_0728_ ) );
INV_X1 \malu/Shift/_1287_ ( .A(\malu/Shift/_0204_ ), .ZN(\malu/Shift/_0521_ ) );
AOI21_X1 \malu/Shift/_1288_ ( .A(\malu/Shift/_0402_ ), .B1(\malu/Shift/_0521_ ), .B2(\malu/Shift/_0720_ ), .ZN(\malu/Shift/_0522_ ) );
OAI21_X1 \malu/Shift/_1289_ ( .A(\malu/Shift/_0034_ ), .B1(\malu/Shift/_0119_ ), .B2(\malu/Shift/_0178_ ), .ZN(\malu/Shift/_0523_ ) );
OAI21_X1 \malu/Shift/_1290_ ( .A(\malu/Shift/_0717_ ), .B1(\malu/Shift/_0176_ ), .B2(\malu/Shift/_0173_ ), .ZN(\malu/Shift/_0524_ ) );
NAND3_X1 \malu/Shift/_1291_ ( .A1(\malu/Shift/_0523_ ), .A2(\malu/Shift/_0052_ ), .A3(\malu/Shift/_0524_ ), .ZN(\malu/Shift/_0525_ ) );
NAND3_X1 \malu/Shift/_1292_ ( .A1(\malu/Shift/_0473_ ), .A2(\malu/Shift/_0474_ ), .A3(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0526_ ) );
AND2_X1 \malu/Shift/_1293_ ( .A1(\malu/Shift/_0525_ ), .A2(\malu/Shift/_0526_ ), .ZN(\malu/Shift/_0527_ ) );
MUX2_X1 \malu/Shift/_1294_ ( .A(\malu/Shift/_0527_ ), .B(\malu/Shift/_0420_ ), .S(\malu/Shift/_0719_ ), .Z(\malu/Shift/_0528_ ) );
OAI21_X1 \malu/Shift/_1295_ ( .A(\malu/Shift/_0522_ ), .B1(\malu/Shift/_0528_ ), .B2(\malu/Shift/_0720_ ), .ZN(\malu/Shift/_0529_ ) );
OR3_X1 \malu/Shift/_1296_ ( .A1(\malu/Shift/_0147_ ), .A2(\malu/Shift/_0720_ ), .A3(\malu/Shift/_0308_ ), .ZN(\malu/Shift/_0530_ ) );
AND2_X1 \malu/Shift/_1297_ ( .A1(\malu/Shift/_0194_ ), .A2(\malu/Shift/_0108_ ), .ZN(\malu/Shift/_0531_ ) );
OAI21_X1 \malu/Shift/_1298_ ( .A(\malu/Shift/_0531_ ), .B1(\malu/Shift/_0200_ ), .B2(\malu/Shift/_0133_ ), .ZN(\malu/Shift/_0532_ ) );
AOI22_X1 \malu/Shift/_1299_ ( .A1(\malu/Shift/_0113_ ), .A2(\malu/Shift/_0507_ ), .B1(\malu/Shift/_0635_ ), .B2(\malu/Shift/_0008_ ), .ZN(\malu/Shift/_0533_ ) );
NAND4_X1 \malu/Shift/_1300_ ( .A1(\malu/Shift/_0529_ ), .A2(\malu/Shift/_0530_ ), .A3(\malu/Shift/_0532_ ), .A4(\malu/Shift/_0533_ ), .ZN(\malu/Shift/_0729_ ) );
OR3_X1 \malu/Shift/_1301_ ( .A1(\malu/Shift/_0224_ ), .A2(\malu/Shift/_0720_ ), .A3(\malu/Shift/_0308_ ), .ZN(\malu/Shift/_0534_ ) );
OAI21_X1 \malu/Shift/_1302_ ( .A(\malu/Shift/_0531_ ), .B1(\malu/Shift/_0216_ ), .B2(\malu/Shift/_0244_ ), .ZN(\malu/Shift/_0535_ ) );
AND3_X2 \malu/Shift/_1303_ ( .A1(\malu/Shift/_0534_ ), .A2(\malu/Shift/_0518_ ), .A3(\malu/Shift/_0535_ ), .ZN(\malu/Shift/_0536_ ) );
NOR4_X1 \malu/Shift/_1304_ ( .A1(\malu/Shift/_0247_ ), .A2(\malu/Shift/_0148_ ), .A3(\malu/Shift/_0718_ ), .A4(\malu/Shift/_0719_ ), .ZN(\malu/Shift/_0537_ ) );
NAND2_X1 \malu/Shift/_1305_ ( .A1(\malu/Shift/_0435_ ), .A2(\malu/Shift/_0438_ ), .ZN(\malu/Shift/_0538_ ) );
OAI21_X1 \malu/Shift/_1306_ ( .A(\malu/Shift/_0717_ ), .B1(\malu/Shift/_0073_ ), .B2(\malu/Shift/_0707_ ), .ZN(\malu/Shift/_0539_ ) );
OAI21_X1 \malu/Shift/_1307_ ( .A(\malu/Shift/_0034_ ), .B1(\malu/Shift/_0077_ ), .B2(\malu/Shift/_0074_ ), .ZN(\malu/Shift/_0540_ ) );
NAND2_X1 \malu/Shift/_1308_ ( .A1(\malu/Shift/_0539_ ), .A2(\malu/Shift/_0540_ ), .ZN(\malu/Shift/_0541_ ) );
NAND2_X1 \malu/Shift/_1309_ ( .A1(\malu/Shift/_0541_ ), .A2(\malu/Shift/_0151_ ), .ZN(\malu/Shift/_0542_ ) );
NAND3_X1 \malu/Shift/_1310_ ( .A1(\malu/Shift/_0487_ ), .A2(\malu/Shift/_0488_ ), .A3(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0543_ ) );
NAND2_X1 \malu/Shift/_1311_ ( .A1(\malu/Shift/_0542_ ), .A2(\malu/Shift/_0543_ ), .ZN(\malu/Shift/_0544_ ) );
MUX2_X1 \malu/Shift/_1312_ ( .A(\malu/Shift/_0538_ ), .B(\malu/Shift/_0544_ ), .S(\malu/Shift/_0236_ ), .Z(\malu/Shift/_0545_ ) );
AOI21_X1 \malu/Shift/_1313_ ( .A(\malu/Shift/_0537_ ), .B1(\malu/Shift/_0545_ ), .B2(\malu/Shift/_0149_ ), .ZN(\malu/Shift/_0546_ ) );
OAI221_X1 \malu/Shift/_1314_ ( .A(\malu/Shift/_0536_ ), .B1(\malu/Shift/_0076_ ), .B2(\malu/Shift/_0104_ ), .C1(\malu/Shift/_0402_ ), .C2(\malu/Shift/_0546_ ), .ZN(\malu/Shift/_0730_ ) );
OR3_X1 \malu/Shift/_1315_ ( .A1(\malu/Shift/_0263_ ), .A2(\malu/Shift/_0720_ ), .A3(\malu/Shift/_0308_ ), .ZN(\malu/Shift/_0547_ ) );
NAND3_X1 \malu/Shift/_1316_ ( .A1(\malu/Shift/_0120_ ), .A2(\malu/Shift/_0717_ ), .A3(\malu/Shift/_0179_ ), .ZN(\malu/Shift/_0548_ ) );
NAND3_X1 \malu/Shift/_1317_ ( .A1(\malu/Shift/_0115_ ), .A2(\malu/Shift/_0038_ ), .A3(\malu/Shift/_0122_ ), .ZN(\malu/Shift/_0549_ ) );
AND2_X1 \malu/Shift/_1318_ ( .A1(\malu/Shift/_0548_ ), .A2(\malu/Shift/_0549_ ), .ZN(\malu/Shift/_0550_ ) );
MUX2_X1 \malu/Shift/_1319_ ( .A(\malu/Shift/_0500_ ), .B(\malu/Shift/_0550_ ), .S(\malu/Shift/_0080_ ), .Z(\malu/Shift/_0551_ ) );
MUX2_X1 \malu/Shift/_1320_ ( .A(\malu/Shift/_0455_ ), .B(\malu/Shift/_0551_ ), .S(\malu/Shift/_0048_ ), .Z(\malu/Shift/_0552_ ) );
NAND2_X1 \malu/Shift/_1321_ ( .A1(\malu/Shift/_0552_ ), .A2(\malu/Shift/_0205_ ), .ZN(\malu/Shift/_0553_ ) );
AND2_X2 \malu/Shift/_1322_ ( .A1(\malu/Shift/_0646_ ), .A2(\malu/Shift/_0720_ ), .ZN(\malu/Shift/_0554_ ) );
AOI221_X4 \malu/Shift/_1323_ ( .A(\malu/Shift/_0517_ ), .B1(\malu/Shift/_0010_ ), .B2(\malu/Shift/_0635_ ), .C1(\malu/Shift/_0290_ ), .C2(\malu/Shift/_0554_ ), .ZN(\malu/Shift/_0555_ ) );
OAI21_X1 \malu/Shift/_1324_ ( .A(\malu/Shift/_0531_ ), .B1(\malu/Shift/_0285_ ), .B2(\malu/Shift/_0262_ ), .ZN(\malu/Shift/_0556_ ) );
NAND4_X1 \malu/Shift/_1325_ ( .A1(\malu/Shift/_0547_ ), .A2(\malu/Shift/_0553_ ), .A3(\malu/Shift/_0555_ ), .A4(\malu/Shift/_0556_ ), .ZN(\malu/Shift/_0731_ ) );
OR2_X1 \malu/Shift/_1326_ ( .A1(\malu/Shift/_0299_ ), .A2(\malu/Shift/_0109_ ), .ZN(\malu/Shift/_0557_ ) );
NAND3_X1 \malu/Shift/_1327_ ( .A1(\malu/Shift/_0510_ ), .A2(\malu/Shift/_0718_ ), .A3(\malu/Shift/_0511_ ), .ZN(\malu/Shift/_0558_ ) );
OR3_X1 \malu/Shift/_1328_ ( .A1(\malu/Shift/_0077_ ), .A2(\malu/Shift/_0074_ ), .A3(\malu/Shift/_0038_ ), .ZN(\malu/Shift/_0559_ ) );
OAI211_X2 \malu/Shift/_1329_ ( .A(\malu/Shift/_0208_ ), .B(\malu/Shift/_0034_ ), .C1(\malu/Shift/_0716_ ), .C2(\malu/Shift/_0068_ ), .ZN(\malu/Shift/_0560_ ) );
NAND3_X1 \malu/Shift/_1330_ ( .A1(\malu/Shift/_0559_ ), .A2(\malu/Shift/_0560_ ), .A3(\malu/Shift/_0151_ ), .ZN(\malu/Shift/_0561_ ) );
NAND2_X1 \malu/Shift/_1331_ ( .A1(\malu/Shift/_0558_ ), .A2(\malu/Shift/_0561_ ), .ZN(\malu/Shift/_0562_ ) );
MUX2_X1 \malu/Shift/_1332_ ( .A(\malu/Shift/_0463_ ), .B(\malu/Shift/_0562_ ), .S(\malu/Shift/_0048_ ), .Z(\malu/Shift/_0563_ ) );
OAI21_X1 \malu/Shift/_1333_ ( .A(\malu/Shift/_0557_ ), .B1(\malu/Shift/_0563_ ), .B2(\malu/Shift/_0720_ ), .ZN(\malu/Shift/_0564_ ) );
OAI21_X1 \malu/Shift/_1334_ ( .A(\malu/Shift/_0149_ ), .B1(\malu/Shift/_0315_ ), .B2(\malu/Shift/_0318_ ), .ZN(\malu/Shift/_0565_ ) );
NAND3_X1 \malu/Shift/_1335_ ( .A1(\malu/Shift/_0714_ ), .A2(\malu/Shift/_0715_ ), .A3(\malu/Shift/_0012_ ), .ZN(\malu/Shift/_0566_ ) );
NAND4_X1 \malu/Shift/_1336_ ( .A1(\malu/Shift/_0564_ ), .A2(\malu/Shift/_0518_ ), .A3(\malu/Shift/_0565_ ), .A4(\malu/Shift/_0566_ ), .ZN(\malu/Shift/_0733_ ) );
AND2_X2 \malu/Shift/_1337_ ( .A1(\malu/Shift/_0328_ ), .A2(\malu/Shift/_0148_ ), .ZN(\malu/Shift/_0567_ ) );
OAI211_X2 \malu/Shift/_1338_ ( .A(\malu/Shift/_0719_ ), .B(\malu/Shift/_0475_ ), .C1(\malu/Shift/_0418_ ), .C2(\malu/Shift/_0053_ ), .ZN(\malu/Shift/_0568_ ) );
OAI21_X1 \malu/Shift/_1339_ ( .A(\malu/Shift/_0034_ ), .B1(\malu/Shift/_0125_ ), .B2(\malu/Shift/_0116_ ), .ZN(\malu/Shift/_0569_ ) );
OAI21_X1 \malu/Shift/_1340_ ( .A(\malu/Shift/_0717_ ), .B1(\malu/Shift/_0114_ ), .B2(\malu/Shift/_0121_ ), .ZN(\malu/Shift/_0570_ ) );
AOI21_X1 \malu/Shift/_1341_ ( .A(\malu/Shift/_0718_ ), .B1(\malu/Shift/_0569_ ), .B2(\malu/Shift/_0570_ ), .ZN(\malu/Shift/_0571_ ) );
AOI21_X1 \malu/Shift/_1342_ ( .A(\malu/Shift/_0052_ ), .B1(\malu/Shift/_0523_ ), .B2(\malu/Shift/_0524_ ), .ZN(\malu/Shift/_0572_ ) );
OAI21_X1 \malu/Shift/_1343_ ( .A(\malu/Shift/_0064_ ), .B1(\malu/Shift/_0571_ ), .B2(\malu/Shift/_0572_ ), .ZN(\malu/Shift/_0573_ ) );
AOI21_X1 \malu/Shift/_1344_ ( .A(\malu/Shift/_0110_ ), .B1(\malu/Shift/_0568_ ), .B2(\malu/Shift/_0573_ ), .ZN(\malu/Shift/_0574_ ) );
AND3_X1 \malu/Shift/_1345_ ( .A1(\malu/Shift/_0345_ ), .A2(\malu/Shift/_0236_ ), .A3(\malu/Shift/_0554_ ), .ZN(\malu/Shift/_0575_ ) );
NAND3_X1 \malu/Shift/_1346_ ( .A1(\malu/Shift/_0714_ ), .A2(\malu/Shift/_0715_ ), .A3(\malu/Shift/_0013_ ), .ZN(\malu/Shift/_0576_ ) );
NAND2_X1 \malu/Shift/_1347_ ( .A1(\malu/Shift/_0112_ ), .A2(\malu/Shift/_0024_ ), .ZN(\malu/Shift/_0577_ ) );
OAI21_X1 \malu/Shift/_1348_ ( .A(\malu/Shift/_0576_ ), .B1(\malu/Shift/_0577_ ), .B2(\malu/Shift/_0148_ ), .ZN(\malu/Shift/_0578_ ) );
OR4_X2 \malu/Shift/_1349_ ( .A1(\malu/Shift/_0567_ ), .A2(\malu/Shift/_0574_ ), .A3(\malu/Shift/_0575_ ), .A4(\malu/Shift/_0578_ ), .ZN(\malu/Shift/_0734_ ) );
NAND2_X1 \malu/Shift/_1350_ ( .A1(\malu/Shift/_0355_ ), .A2(\malu/Shift/_0149_ ), .ZN(\malu/Shift/_0579_ ) );
AOI221_X4 \malu/Shift/_1351_ ( .A(\malu/Shift/_0517_ ), .B1(\malu/Shift/_0014_ ), .B2(\malu/Shift/_0635_ ), .C1(\malu/Shift/_0368_ ), .C2(\malu/Shift/_0554_ ), .ZN(\malu/Shift/_0580_ ) );
NAND2_X1 \malu/Shift/_1352_ ( .A1(\malu/Shift/_0541_ ), .A2(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0581_ ) );
OR3_X1 \malu/Shift/_1353_ ( .A1(\malu/Shift/_0065_ ), .A2(\malu/Shift/_0070_ ), .A3(\malu/Shift/_0717_ ), .ZN(\malu/Shift/_0582_ ) );
OAI211_X2 \malu/Shift/_1354_ ( .A(\malu/Shift/_0208_ ), .B(\malu/Shift/_0717_ ), .C1(\malu/Shift/_0716_ ), .C2(\malu/Shift/_0068_ ), .ZN(\malu/Shift/_0583_ ) );
NAND3_X1 \malu/Shift/_1355_ ( .A1(\malu/Shift/_0582_ ), .A2(\malu/Shift/_0583_ ), .A3(\malu/Shift/_0052_ ), .ZN(\malu/Shift/_0584_ ) );
AOI21_X1 \malu/Shift/_1356_ ( .A(\malu/Shift/_0719_ ), .B1(\malu/Shift/_0581_ ), .B2(\malu/Shift/_0584_ ), .ZN(\malu/Shift/_0585_ ) );
AOI21_X1 \malu/Shift/_1357_ ( .A(\malu/Shift/_0585_ ), .B1(\malu/Shift/_0719_ ), .B2(\malu/Shift/_0490_ ), .ZN(\malu/Shift/_0586_ ) );
OAI211_X2 \malu/Shift/_1358_ ( .A(\malu/Shift/_0579_ ), .B(\malu/Shift/_0580_ ), .C1(\malu/Shift/_0110_ ), .C2(\malu/Shift/_0586_ ), .ZN(\malu/Shift/_0735_ ) );
AOI21_X1 \malu/Shift/_1359_ ( .A(\malu/Shift/_0151_ ), .B1(\malu/Shift/_0548_ ), .B2(\malu/Shift/_0549_ ), .ZN(\malu/Shift/_0587_ ) );
OAI21_X1 \malu/Shift/_1360_ ( .A(\malu/Shift/_0034_ ), .B1(\malu/Shift/_0128_ ), .B2(\malu/Shift/_0126_ ), .ZN(\malu/Shift/_0588_ ) );
OAI21_X1 \malu/Shift/_1361_ ( .A(\malu/Shift/_0717_ ), .B1(\malu/Shift/_0125_ ), .B2(\malu/Shift/_0116_ ), .ZN(\malu/Shift/_0589_ ) );
AND3_X1 \malu/Shift/_1362_ ( .A1(\malu/Shift/_0588_ ), .A2(\malu/Shift/_0589_ ), .A3(\malu/Shift/_0052_ ), .ZN(\malu/Shift/_0590_ ) );
OAI21_X1 \malu/Shift/_1363_ ( .A(\malu/Shift/_0236_ ), .B1(\malu/Shift/_0587_ ), .B2(\malu/Shift/_0590_ ), .ZN(\malu/Shift/_0591_ ) );
NAND3_X1 \malu/Shift/_1364_ ( .A1(\malu/Shift/_0501_ ), .A2(\malu/Shift/_0502_ ), .A3(\malu/Shift/_0719_ ), .ZN(\malu/Shift/_0592_ ) );
AND3_X1 \malu/Shift/_1365_ ( .A1(\malu/Shift/_0591_ ), .A2(\malu/Shift/_0249_ ), .A3(\malu/Shift/_0592_ ), .ZN(\malu/Shift/_0593_ ) );
OAI21_X1 \malu/Shift/_1366_ ( .A(\malu/Shift/_0149_ ), .B1(\malu/Shift/_0377_ ), .B2(\malu/Shift/_0593_ ), .ZN(\malu/Shift/_0594_ ) );
NAND3_X1 \malu/Shift/_1367_ ( .A1(\malu/Shift/_0390_ ), .A2(\malu/Shift/_0335_ ), .A3(\malu/Shift/_0554_ ), .ZN(\malu/Shift/_0595_ ) );
NAND3_X1 \malu/Shift/_1368_ ( .A1(\malu/Shift/_0714_ ), .A2(\malu/Shift/_0715_ ), .A3(\malu/Shift/_0015_ ), .ZN(\malu/Shift/_0596_ ) );
NAND4_X1 \malu/Shift/_1369_ ( .A1(\malu/Shift/_0594_ ), .A2(\malu/Shift/_0518_ ), .A3(\malu/Shift/_0595_ ), .A4(\malu/Shift/_0596_ ), .ZN(\malu/Shift/_0736_ ) );
NAND3_X1 \malu/Shift/_1370_ ( .A1(\malu/Shift/_0395_ ), .A2(\malu/Shift/_0397_ ), .A3(\malu/Shift/_0518_ ), .ZN(\malu/Shift/_0597_ ) );
NAND2_X1 \malu/Shift/_1371_ ( .A1(\malu/Shift/_0577_ ), .A2(\malu/Shift/_0720_ ), .ZN(\malu/Shift/_0598_ ) );
NAND2_X1 \malu/Shift/_1372_ ( .A1(\malu/Shift/_0597_ ), .A2(\malu/Shift/_0598_ ), .ZN(\malu/Shift/_0599_ ) );
NAND2_X1 \malu/Shift/_1373_ ( .A1(\malu/Shift/_0410_ ), .A2(\malu/Shift/_0110_ ), .ZN(\malu/Shift/_0600_ ) );
OR3_X1 \malu/Shift/_1374_ ( .A1(\malu/Shift/_0065_ ), .A2(\malu/Shift/_0070_ ), .A3(\malu/Shift/_0038_ ), .ZN(\malu/Shift/_0601_ ) );
NOR2_X1 \malu/Shift/_1375_ ( .A1(\malu/Shift/_0085_ ), .A2(\malu/Shift/_0716_ ), .ZN(\malu/Shift/_0602_ ) );
OR3_X1 \malu/Shift/_1376_ ( .A1(\malu/Shift/_0602_ ), .A2(\malu/Shift/_0066_ ), .A3(\malu/Shift/_0717_ ), .ZN(\malu/Shift/_0603_ ) );
AOI21_X1 \malu/Shift/_1377_ ( .A(\malu/Shift/_0718_ ), .B1(\malu/Shift/_0601_ ), .B2(\malu/Shift/_0603_ ), .ZN(\malu/Shift/_0604_ ) );
AOI21_X1 \malu/Shift/_1378_ ( .A(\malu/Shift/_0052_ ), .B1(\malu/Shift/_0559_ ), .B2(\malu/Shift/_0560_ ), .ZN(\malu/Shift/_0605_ ) );
NOR2_X1 \malu/Shift/_1379_ ( .A1(\malu/Shift/_0604_ ), .A2(\malu/Shift/_0605_ ), .ZN(\malu/Shift/_0606_ ) );
MUX2_X1 \malu/Shift/_1380_ ( .A(\malu/Shift/_0514_ ), .B(\malu/Shift/_0606_ ), .S(\malu/Shift/_0064_ ), .Z(\malu/Shift/_0607_ ) );
OAI21_X1 \malu/Shift/_1381_ ( .A(\malu/Shift/_0600_ ), .B1(\malu/Shift/_0607_ ), .B2(\malu/Shift/_0720_ ), .ZN(\malu/Shift/_0608_ ) );
OAI211_X2 \malu/Shift/_1382_ ( .A(\malu/Shift/_0599_ ), .B(\malu/Shift/_0608_ ), .C1(\malu/Shift/_0085_ ), .C2(\malu/Shift/_0105_ ), .ZN(\malu/Shift/_0737_ ) );
NAND2_X1 \malu/Shift/_1383_ ( .A1(\malu/Shift/_0421_ ), .A2(\malu/Shift/_0249_ ), .ZN(\malu/Shift/_0609_ ) );
NAND2_X1 \malu/Shift/_1384_ ( .A1(\malu/Shift/_0609_ ), .A2(\malu/Shift/_0110_ ), .ZN(\malu/Shift/_0610_ ) );
AND3_X1 \malu/Shift/_1385_ ( .A1(\malu/Shift/_0569_ ), .A2(\malu/Shift/_0570_ ), .A3(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0611_ ) );
OR3_X1 \malu/Shift/_1386_ ( .A1(\malu/Shift/_0128_ ), .A2(\malu/Shift/_0033_ ), .A3(\malu/Shift/_0126_ ), .ZN(\malu/Shift/_0612_ ) );
OR3_X1 \malu/Shift/_1387_ ( .A1(\malu/Shift/_0139_ ), .A2(\malu/Shift/_0717_ ), .A3(\malu/Shift/_0129_ ), .ZN(\malu/Shift/_0613_ ) );
AND2_X1 \malu/Shift/_1388_ ( .A1(\malu/Shift/_0612_ ), .A2(\malu/Shift/_0613_ ), .ZN(\malu/Shift/_0614_ ) );
INV_X1 \malu/Shift/_1389_ ( .A(\malu/Shift/_0614_ ), .ZN(\malu/Shift/_0615_ ) );
AOI21_X1 \malu/Shift/_1390_ ( .A(\malu/Shift/_0611_ ), .B1(\malu/Shift/_0615_ ), .B2(\malu/Shift/_0100_ ), .ZN(\malu/Shift/_0616_ ) );
MUX2_X1 \malu/Shift/_1391_ ( .A(\malu/Shift/_0527_ ), .B(\malu/Shift/_0616_ ), .S(\malu/Shift/_0236_ ), .Z(\malu/Shift/_0617_ ) );
OAI21_X1 \malu/Shift/_1392_ ( .A(\malu/Shift/_0610_ ), .B1(\malu/Shift/_0720_ ), .B2(\malu/Shift/_0617_ ), .ZN(\malu/Shift/_0618_ ) );
AOI21_X1 \malu/Shift/_1393_ ( .A(\malu/Shift/_0720_ ), .B1(\malu/Shift/_0423_ ), .B2(\malu/Shift/_0424_ ), .ZN(\malu/Shift/_0619_ ) );
OAI21_X1 \malu/Shift/_1394_ ( .A(\malu/Shift/_0113_ ), .B1(\malu/Shift/_0619_ ), .B2(\malu/Shift/_0507_ ), .ZN(\malu/Shift/_0620_ ) );
OR4_X4 \malu/Shift/_1395_ ( .A1(\malu/Shift/_0720_ ), .A2(\malu/Shift/_0199_ ), .A3(\malu/Shift/_0719_ ), .A4(\malu/Shift/_0316_ ), .ZN(\malu/Shift/_0621_ ) );
NAND3_X1 \malu/Shift/_1396_ ( .A1(\malu/Shift/_0714_ ), .A2(\malu/Shift/_0715_ ), .A3(\malu/Shift/_0017_ ), .ZN(\malu/Shift/_0622_ ) );
NAND4_X1 \malu/Shift/_1397_ ( .A1(\malu/Shift/_0618_ ), .A2(\malu/Shift/_0620_ ), .A3(\malu/Shift/_0621_ ), .A4(\malu/Shift/_0622_ ), .ZN(\malu/Shift/_0738_ ) );
OAI211_X2 \malu/Shift/_1398_ ( .A(\malu/Shift/_0432_ ), .B(\malu/Shift/_0518_ ), .C1(\malu/Shift/_0308_ ), .C2(\malu/Shift/_0429_ ), .ZN(\malu/Shift/_0623_ ) );
NAND2_X1 \malu/Shift/_1399_ ( .A1(\malu/Shift/_0623_ ), .A2(\malu/Shift/_0598_ ), .ZN(\malu/Shift/_0624_ ) );
NAND3_X1 \malu/Shift/_1400_ ( .A1(\malu/Shift/_0582_ ), .A2(\malu/Shift/_0583_ ), .A3(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0625_ ) );
NOR2_X1 \malu/Shift/_1401_ ( .A1(\malu/Shift/_0217_ ), .A2(\malu/Shift/_0083_ ), .ZN(\malu/Shift/_0626_ ) );
NOR2_X1 \malu/Shift/_1402_ ( .A1(\malu/Shift/_0602_ ), .A2(\malu/Shift/_0066_ ), .ZN(\malu/Shift/_0627_ ) );
MUX2_X1 \malu/Shift/_1403_ ( .A(\malu/Shift/_0626_ ), .B(\malu/Shift/_0627_ ), .S(\malu/Shift/_0717_ ), .Z(\malu/Shift/_0628_ ) );
OAI211_X2 \malu/Shift/_1404_ ( .A(\malu/Shift/_0625_ ), .B(\malu/Shift/_0236_ ), .C1(\malu/Shift/_0628_ ), .C2(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0629_ ) );
AND2_X1 \malu/Shift/_1405_ ( .A1(\malu/Shift/_0629_ ), .A2(\malu/Shift/_0205_ ), .ZN(\malu/Shift/_0630_ ) );
OAI21_X1 \malu/Shift/_1406_ ( .A(\malu/Shift/_0630_ ), .B1(\malu/Shift/_0335_ ), .B2(\malu/Shift/_0544_ ), .ZN(\malu/Shift/_0631_ ) );
NAND3_X1 \malu/Shift/_1407_ ( .A1(\malu/Shift/_0714_ ), .A2(\malu/Shift/_0715_ ), .A3(\malu/Shift/_0018_ ), .ZN(\malu/Shift/_0632_ ) );
OAI21_X1 \malu/Shift/_1408_ ( .A(\malu/Shift/_0554_ ), .B1(\malu/Shift/_0434_ ), .B2(\malu/Shift/_0439_ ), .ZN(\malu/Shift/_0633_ ) );
NAND4_X1 \malu/Shift/_1409_ ( .A1(\malu/Shift/_0624_ ), .A2(\malu/Shift/_0631_ ), .A3(\malu/Shift/_0632_ ), .A4(\malu/Shift/_0633_ ), .ZN(\malu/Shift/_0739_ ) );
NAND3_X1 \malu/Shift/_1410_ ( .A1(\malu/Shift/_0444_ ), .A2(\malu/Shift/_0445_ ), .A3(\malu/Shift/_0518_ ), .ZN(\malu/Shift/_0634_ ) );
AND2_X1 \malu/Shift/_1411_ ( .A1(\malu/Shift/_0634_ ), .A2(\malu/Shift/_0598_ ), .ZN(\malu/Shift/_0636_ ) );
NAND2_X1 \malu/Shift/_1412_ ( .A1(\malu/Shift/_0551_ ), .A2(\malu/Shift/_0719_ ), .ZN(\malu/Shift/_0637_ ) );
NAND3_X1 \malu/Shift/_1413_ ( .A1(\malu/Shift/_0588_ ), .A2(\malu/Shift/_0589_ ), .A3(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0638_ ) );
OAI21_X1 \malu/Shift/_1414_ ( .A(\malu/Shift/_0039_ ), .B1(\malu/Shift/_0142_ ), .B2(\malu/Shift/_0140_ ), .ZN(\malu/Shift/_0639_ ) );
OAI21_X1 \malu/Shift/_1415_ ( .A(\malu/Shift/_0717_ ), .B1(\malu/Shift/_0139_ ), .B2(\malu/Shift/_0129_ ), .ZN(\malu/Shift/_0640_ ) );
NAND2_X1 \malu/Shift/_1416_ ( .A1(\malu/Shift/_0639_ ), .A2(\malu/Shift/_0640_ ), .ZN(\malu/Shift/_0641_ ) );
OAI211_X2 \malu/Shift/_1417_ ( .A(\malu/Shift/_0638_ ), .B(\malu/Shift/_0064_ ), .C1(\malu/Shift/_0641_ ), .C2(\malu/Shift/_0718_ ), .ZN(\malu/Shift/_0642_ ) );
AOI21_X1 \malu/Shift/_1418_ ( .A(\malu/Shift/_0110_ ), .B1(\malu/Shift/_0637_ ), .B2(\malu/Shift/_0642_ ), .ZN(\malu/Shift/_0643_ ) );
AND3_X1 \malu/Shift/_1419_ ( .A1(\malu/Shift/_0714_ ), .A2(\malu/Shift/_0715_ ), .A3(\malu/Shift/_0019_ ), .ZN(\malu/Shift/_0644_ ) );
AND2_X1 \malu/Shift/_1420_ ( .A1(\malu/Shift/_0457_ ), .A2(\malu/Shift/_0554_ ), .ZN(\malu/Shift/_0645_ ) );
OR4_X1 \malu/Shift/_1421_ ( .A1(\malu/Shift/_0636_ ), .A2(\malu/Shift/_0643_ ), .A3(\malu/Shift/_0644_ ), .A4(\malu/Shift/_0645_ ), .ZN(\malu/Shift/_0740_ ) );
AND2_X1 \malu/Shift/_1422_ ( .A1(\malu/Shift/_0468_ ), .A2(\malu/Shift/_0113_ ), .ZN(\malu/Shift/_0647_ ) );
NAND2_X1 \malu/Shift/_1423_ ( .A1(\malu/Shift/_0309_ ), .A2(\malu/Shift/_0396_ ), .ZN(\malu/Shift/_0648_ ) );
NAND2_X1 \malu/Shift/_1424_ ( .A1(\malu/Shift/_0648_ ), .A2(\malu/Shift/_0518_ ), .ZN(\malu/Shift/_0649_ ) );
OAI21_X1 \malu/Shift/_1425_ ( .A(\malu/Shift/_0598_ ), .B1(\malu/Shift/_0647_ ), .B2(\malu/Shift/_0649_ ), .ZN(\malu/Shift/_0650_ ) );
NAND3_X1 \malu/Shift/_1426_ ( .A1(\malu/Shift/_0464_ ), .A2(\malu/Shift/_0720_ ), .A3(\malu/Shift/_0249_ ), .ZN(\malu/Shift/_0651_ ) );
NAND3_X1 \malu/Shift/_1427_ ( .A1(\malu/Shift/_0714_ ), .A2(\malu/Shift/_0715_ ), .A3(\malu/Shift/_0020_ ), .ZN(\malu/Shift/_0652_ ) );
AOI21_X1 \malu/Shift/_1428_ ( .A(\malu/Shift/_0100_ ), .B1(\malu/Shift/_0601_ ), .B2(\malu/Shift/_0603_ ), .ZN(\malu/Shift/_0653_ ) );
OAI211_X2 \malu/Shift/_1429_ ( .A(\malu/Shift/_0088_ ), .B(\malu/Shift/_0039_ ), .C1(\malu/Shift/_0716_ ), .C2(\malu/Shift/_0092_ ), .ZN(\malu/Shift/_0654_ ) );
OAI211_X2 \malu/Shift/_1430_ ( .A(\malu/Shift/_0084_ ), .B(\malu/Shift/_0717_ ), .C1(\malu/Shift/_0716_ ), .C2(\malu/Shift/_0089_ ), .ZN(\malu/Shift/_0655_ ) );
AOI21_X1 \malu/Shift/_1431_ ( .A(\malu/Shift/_0718_ ), .B1(\malu/Shift/_0654_ ), .B2(\malu/Shift/_0655_ ), .ZN(\malu/Shift/_0657_ ) );
OAI21_X1 \malu/Shift/_1432_ ( .A(\malu/Shift/_0236_ ), .B1(\malu/Shift/_0653_ ), .B2(\malu/Shift/_0657_ ), .ZN(\malu/Shift/_0658_ ) );
AND2_X1 \malu/Shift/_1433_ ( .A1(\malu/Shift/_0658_ ), .A2(\malu/Shift/_0109_ ), .ZN(\malu/Shift/_0659_ ) );
OAI21_X1 \malu/Shift/_1434_ ( .A(\malu/Shift/_0659_ ), .B1(\malu/Shift/_0335_ ), .B2(\malu/Shift/_0562_ ), .ZN(\malu/Shift/_0660_ ) );
NAND4_X1 \malu/Shift/_1435_ ( .A1(\malu/Shift/_0650_ ), .A2(\malu/Shift/_0651_ ), .A3(\malu/Shift/_0652_ ), .A4(\malu/Shift/_0660_ ), .ZN(\malu/Shift/_0741_ ) );
OAI21_X1 \malu/Shift/_1436_ ( .A(\malu/Shift/_0598_ ), .B1(\malu/Shift/_0482_ ), .B2(\malu/Shift/_0517_ ), .ZN(\malu/Shift/_0661_ ) );
OR3_X1 \malu/Shift/_1437_ ( .A1(\malu/Shift/_0142_ ), .A2(\malu/Shift/_0039_ ), .A3(\malu/Shift/_0140_ ), .ZN(\malu/Shift/_0662_ ) );
MUX2_X1 \malu/Shift/_1438_ ( .A(\malu/Shift/_0021_ ), .B(\malu/Shift/_0020_ ), .S(\malu/Shift/_0716_ ), .Z(\malu/Shift/_0663_ ) );
OAI211_X2 \malu/Shift/_1439_ ( .A(\malu/Shift/_0662_ ), .B(\malu/Shift/_0053_ ), .C1(\malu/Shift/_0717_ ), .C2(\malu/Shift/_0663_ ), .ZN(\malu/Shift/_0664_ ) );
OAI211_X2 \malu/Shift/_1440_ ( .A(\malu/Shift/_0335_ ), .B(\malu/Shift/_0664_ ), .C1(\malu/Shift/_0615_ ), .C2(\malu/Shift/_0053_ ), .ZN(\malu/Shift/_0665_ ) );
OR3_X1 \malu/Shift/_1441_ ( .A1(\malu/Shift/_0571_ ), .A2(\malu/Shift/_0572_ ), .A3(\malu/Shift/_0236_ ), .ZN(\malu/Shift/_0667_ ) );
NAND3_X1 \malu/Shift/_1442_ ( .A1(\malu/Shift/_0665_ ), .A2(\malu/Shift/_0205_ ), .A3(\malu/Shift/_0667_ ), .ZN(\malu/Shift/_0668_ ) );
NAND3_X1 \malu/Shift/_1443_ ( .A1(\malu/Shift/_0714_ ), .A2(\malu/Shift/_0715_ ), .A3(\malu/Shift/_0021_ ), .ZN(\malu/Shift/_0669_ ) );
NAND2_X1 \malu/Shift/_1444_ ( .A1(\malu/Shift/_0477_ ), .A2(\malu/Shift/_0554_ ), .ZN(\malu/Shift/_0670_ ) );
NAND4_X1 \malu/Shift/_1445_ ( .A1(\malu/Shift/_0661_ ), .A2(\malu/Shift/_0668_ ), .A3(\malu/Shift/_0669_ ), .A4(\malu/Shift/_0670_ ), .ZN(\malu/Shift/_0742_ ) );
AOI221_X1 \malu/Shift/_1446_ ( .A(\malu/Shift/_0517_ ), .B1(\malu/Shift/_0352_ ), .B2(\malu/Shift/_0396_ ), .C1(\malu/Shift/_0493_ ), .C2(\malu/Shift/_0112_ ), .ZN(\malu/Shift/_0671_ ) );
AOI21_X1 \malu/Shift/_1447_ ( .A(\malu/Shift/_0671_ ), .B1(\malu/Shift/_0720_ ), .B2(\malu/Shift/_0577_ ), .ZN(\malu/Shift/_0672_ ) );
AND3_X1 \malu/Shift/_1448_ ( .A1(\malu/Shift/_0491_ ), .A2(\malu/Shift/_0720_ ), .A3(\malu/Shift/_0249_ ), .ZN(\malu/Shift/_0673_ ) );
OAI211_X2 \malu/Shift/_1449_ ( .A(\malu/Shift/_0088_ ), .B(\malu/Shift/_0717_ ), .C1(\malu/Shift/_0716_ ), .C2(\malu/Shift/_0092_ ), .ZN(\malu/Shift/_0674_ ) );
MUX2_X1 \malu/Shift/_1450_ ( .A(\malu/Shift/_0023_ ), .B(\malu/Shift/_0021_ ), .S(\malu/Shift/_0716_ ), .Z(\malu/Shift/_0675_ ) );
OAI211_X2 \malu/Shift/_1451_ ( .A(\malu/Shift/_0674_ ), .B(\malu/Shift/_0052_ ), .C1(\malu/Shift/_0717_ ), .C2(\malu/Shift/_0675_ ), .ZN(\malu/Shift/_0677_ ) );
OAI211_X2 \malu/Shift/_1452_ ( .A(\malu/Shift/_0677_ ), .B(\malu/Shift/_0064_ ), .C1(\malu/Shift/_0628_ ), .C2(\malu/Shift/_0100_ ), .ZN(\malu/Shift/_0678_ ) );
NAND3_X1 \malu/Shift/_1453_ ( .A1(\malu/Shift/_0581_ ), .A2(\malu/Shift/_0584_ ), .A3(\malu/Shift/_0719_ ), .ZN(\malu/Shift/_0679_ ) );
NAND3_X1 \malu/Shift/_1454_ ( .A1(\malu/Shift/_0678_ ), .A2(\malu/Shift/_0108_ ), .A3(\malu/Shift/_0679_ ), .ZN(\malu/Shift/_0680_ ) );
OAI22_X1 \malu/Shift/_1455_ ( .A1(\malu/Shift/_0680_ ), .A2(\malu/Shift/_0402_ ), .B1(\malu/Shift/_0096_ ), .B2(\malu/Shift/_0104_ ), .ZN(\malu/Shift/_0681_ ) );
OR3_X1 \malu/Shift/_1456_ ( .A1(\malu/Shift/_0672_ ), .A2(\malu/Shift/_0673_ ), .A3(\malu/Shift/_0681_ ), .ZN(\malu/Shift/_0744_ ) );
MUX2_X1 \malu/Shift/_1457_ ( .A(\malu/Shift/_0024_ ), .B(\malu/Shift/_0023_ ), .S(\malu/Shift/_0716_ ), .Z(\malu/Shift/_0682_ ) );
MUX2_X1 \malu/Shift/_1458_ ( .A(\malu/Shift/_0682_ ), .B(\malu/Shift/_0663_ ), .S(\malu/Shift/_0717_ ), .Z(\malu/Shift/_0683_ ) );
MUX2_X1 \malu/Shift/_1459_ ( .A(\malu/Shift/_0641_ ), .B(\malu/Shift/_0683_ ), .S(\malu/Shift/_0100_ ), .Z(\malu/Shift/_0684_ ) );
OR2_X1 \malu/Shift/_1460_ ( .A1(\malu/Shift/_0684_ ), .A2(\malu/Shift/_0719_ ), .ZN(\malu/Shift/_0685_ ) );
OAI21_X1 \malu/Shift/_1461_ ( .A(\malu/Shift/_0719_ ), .B1(\malu/Shift/_0587_ ), .B2(\malu/Shift/_0590_ ), .ZN(\malu/Shift/_0687_ ) );
NAND3_X1 \malu/Shift/_1462_ ( .A1(\malu/Shift/_0685_ ), .A2(\malu/Shift/_0205_ ), .A3(\malu/Shift/_0687_ ), .ZN(\malu/Shift/_0688_ ) );
NAND3_X1 \malu/Shift/_1463_ ( .A1(\malu/Shift/_0497_ ), .A2(\malu/Shift/_0503_ ), .A3(\malu/Shift/_0554_ ), .ZN(\malu/Shift/_0689_ ) );
NAND3_X1 \malu/Shift/_1464_ ( .A1(\malu/Shift/_0531_ ), .A2(\malu/Shift/_0505_ ), .A3(\malu/Shift/_0335_ ), .ZN(\malu/Shift/_0690_ ) );
NAND2_X1 \malu/Shift/_1465_ ( .A1(\malu/Shift/_0714_ ), .A2(\malu/Shift/_0024_ ), .ZN(\malu/Shift/_0691_ ) );
NAND4_X1 \malu/Shift/_1466_ ( .A1(\malu/Shift/_0688_ ), .A2(\malu/Shift/_0689_ ), .A3(\malu/Shift/_0690_ ), .A4(\malu/Shift/_0691_ ), .ZN(\malu/Shift/_0745_ ) );
BUF_X1 \malu/Shift/_1467_ ( .A(\malu/shift_ctl[0] ), .Z(\malu/Shift/_0714_ ) );
BUF_X1 \malu/Shift/_1468_ ( .A(\malu/shift_ctl[1] ), .Z(\malu/Shift/_0715_ ) );
BUF_X1 \malu/Shift/_1469_ ( .A(\alu_b[4] ), .Z(\malu/Shift/_0720_ ) );
BUF_X1 \malu/Shift/_1470_ ( .A(\alu_b[2] ), .Z(\malu/Shift/_0718_ ) );
BUF_X1 \malu/Shift/_1471_ ( .A(\alu_b[1] ), .Z(\malu/Shift/_0717_ ) );
BUF_X1 \malu/Shift/_1472_ ( .A(\alu_a[0] ), .Z(\malu/Shift/_0000_ ) );
BUF_X1 \malu/Shift/_1473_ ( .A(\alu_a[1] ), .Z(\malu/Shift/_0011_ ) );
BUF_X1 \malu/Shift/_1474_ ( .A(\alu_b[0] ), .Z(\malu/Shift/_0716_ ) );
BUF_X1 \malu/Shift/_1475_ ( .A(\alu_a[2] ), .Z(\malu/Shift/_0022_ ) );
BUF_X1 \malu/Shift/_1476_ ( .A(\alu_a[3] ), .Z(\malu/Shift/_0025_ ) );
BUF_X1 \malu/Shift/_1477_ ( .A(\alu_a[4] ), .Z(\malu/Shift/_0026_ ) );
BUF_X1 \malu/Shift/_1478_ ( .A(\alu_a[5] ), .Z(\malu/Shift/_0027_ ) );
BUF_X1 \malu/Shift/_1479_ ( .A(\alu_a[6] ), .Z(\malu/Shift/_0028_ ) );
BUF_X1 \malu/Shift/_1480_ ( .A(\alu_a[7] ), .Z(\malu/Shift/_0029_ ) );
BUF_X1 \malu/Shift/_1481_ ( .A(\alu_a[8] ), .Z(\malu/Shift/_0030_ ) );
BUF_X1 \malu/Shift/_1482_ ( .A(\alu_a[9] ), .Z(\malu/Shift/_0031_ ) );
BUF_X1 \malu/Shift/_1483_ ( .A(\alu_a[10] ), .Z(\malu/Shift/_0001_ ) );
BUF_X1 \malu/Shift/_1484_ ( .A(\alu_a[11] ), .Z(\malu/Shift/_0002_ ) );
BUF_X1 \malu/Shift/_1485_ ( .A(\alu_a[12] ), .Z(\malu/Shift/_0003_ ) );
BUF_X1 \malu/Shift/_1486_ ( .A(\alu_a[13] ), .Z(\malu/Shift/_0004_ ) );
BUF_X1 \malu/Shift/_1487_ ( .A(\alu_a[14] ), .Z(\malu/Shift/_0005_ ) );
BUF_X1 \malu/Shift/_1488_ ( .A(\alu_a[15] ), .Z(\malu/Shift/_0006_ ) );
BUF_X1 \malu/Shift/_1489_ ( .A(\alu_b[3] ), .Z(\malu/Shift/_0719_ ) );
BUF_X1 \malu/Shift/_1490_ ( .A(\alu_a[16] ), .Z(\malu/Shift/_0007_ ) );
BUF_X1 \malu/Shift/_1491_ ( .A(\alu_a[17] ), .Z(\malu/Shift/_0008_ ) );
BUF_X1 \malu/Shift/_1492_ ( .A(\alu_a[18] ), .Z(\malu/Shift/_0009_ ) );
BUF_X1 \malu/Shift/_1493_ ( .A(\alu_a[19] ), .Z(\malu/Shift/_0010_ ) );
BUF_X1 \malu/Shift/_1494_ ( .A(\alu_a[20] ), .Z(\malu/Shift/_0012_ ) );
BUF_X1 \malu/Shift/_1495_ ( .A(\alu_a[21] ), .Z(\malu/Shift/_0013_ ) );
BUF_X1 \malu/Shift/_1496_ ( .A(\alu_a[22] ), .Z(\malu/Shift/_0014_ ) );
BUF_X1 \malu/Shift/_1497_ ( .A(\alu_a[23] ), .Z(\malu/Shift/_0015_ ) );
BUF_X1 \malu/Shift/_1498_ ( .A(\alu_a[24] ), .Z(\malu/Shift/_0016_ ) );
BUF_X1 \malu/Shift/_1499_ ( .A(\alu_a[25] ), .Z(\malu/Shift/_0017_ ) );
BUF_X1 \malu/Shift/_1500_ ( .A(\alu_a[26] ), .Z(\malu/Shift/_0018_ ) );
BUF_X1 \malu/Shift/_1501_ ( .A(\alu_a[27] ), .Z(\malu/Shift/_0019_ ) );
BUF_X1 \malu/Shift/_1502_ ( .A(\alu_a[28] ), .Z(\malu/Shift/_0020_ ) );
BUF_X1 \malu/Shift/_1503_ ( .A(\alu_a[29] ), .Z(\malu/Shift/_0021_ ) );
BUF_X1 \malu/Shift/_1504_ ( .A(\alu_a[30] ), .Z(\malu/Shift/_0023_ ) );
BUF_X1 \malu/Shift/_1505_ ( .A(\alu_a[31] ), .Z(\malu/Shift/_0024_ ) );
BUF_X1 \malu/Shift/_1506_ ( .A(\malu/Shift/_0721_ ), .Z(\malu/shift_result[0] ) );
BUF_X1 \malu/Shift/_1507_ ( .A(\malu/Shift/_0732_ ), .Z(\malu/shift_result[1] ) );
BUF_X1 \malu/Shift/_1508_ ( .A(\malu/Shift/_0743_ ), .Z(\malu/shift_result[2] ) );
BUF_X1 \malu/Shift/_1509_ ( .A(\malu/Shift/_0746_ ), .Z(\malu/shift_result[3] ) );
BUF_X1 \malu/Shift/_1510_ ( .A(\malu/Shift/_0747_ ), .Z(\malu/shift_result[4] ) );
BUF_X1 \malu/Shift/_1511_ ( .A(\malu/Shift/_0748_ ), .Z(\malu/shift_result[5] ) );
BUF_X1 \malu/Shift/_1512_ ( .A(\malu/Shift/_0749_ ), .Z(\malu/shift_result[6] ) );
BUF_X1 \malu/Shift/_1513_ ( .A(\malu/Shift/_0750_ ), .Z(\malu/shift_result[7] ) );
BUF_X1 \malu/Shift/_1514_ ( .A(\malu/Shift/_0751_ ), .Z(\malu/shift_result[8] ) );
BUF_X1 \malu/Shift/_1515_ ( .A(\malu/Shift/_0752_ ), .Z(\malu/shift_result[9] ) );
BUF_X1 \malu/Shift/_1516_ ( .A(\malu/Shift/_0722_ ), .Z(\malu/shift_result[10] ) );
BUF_X1 \malu/Shift/_1517_ ( .A(\malu/Shift/_0723_ ), .Z(\malu/shift_result[11] ) );
BUF_X1 \malu/Shift/_1518_ ( .A(\malu/Shift/_0724_ ), .Z(\malu/shift_result[12] ) );
BUF_X1 \malu/Shift/_1519_ ( .A(\malu/Shift/_0725_ ), .Z(\malu/shift_result[13] ) );
BUF_X1 \malu/Shift/_1520_ ( .A(\malu/Shift/_0726_ ), .Z(\malu/shift_result[14] ) );
BUF_X1 \malu/Shift/_1521_ ( .A(\malu/Shift/_0727_ ), .Z(\malu/shift_result[15] ) );
BUF_X1 \malu/Shift/_1522_ ( .A(\malu/Shift/_0728_ ), .Z(\malu/shift_result[16] ) );
BUF_X1 \malu/Shift/_1523_ ( .A(\malu/Shift/_0729_ ), .Z(\malu/shift_result[17] ) );
BUF_X1 \malu/Shift/_1524_ ( .A(\malu/Shift/_0730_ ), .Z(\malu/shift_result[18] ) );
BUF_X1 \malu/Shift/_1525_ ( .A(\malu/Shift/_0731_ ), .Z(\malu/shift_result[19] ) );
BUF_X1 \malu/Shift/_1526_ ( .A(\malu/Shift/_0733_ ), .Z(\malu/shift_result[20] ) );
BUF_X1 \malu/Shift/_1527_ ( .A(\malu/Shift/_0734_ ), .Z(\malu/shift_result[21] ) );
BUF_X1 \malu/Shift/_1528_ ( .A(\malu/Shift/_0735_ ), .Z(\malu/shift_result[22] ) );
BUF_X1 \malu/Shift/_1529_ ( .A(\malu/Shift/_0736_ ), .Z(\malu/shift_result[23] ) );
BUF_X1 \malu/Shift/_1530_ ( .A(\malu/Shift/_0737_ ), .Z(\malu/shift_result[24] ) );
BUF_X1 \malu/Shift/_1531_ ( .A(\malu/Shift/_0738_ ), .Z(\malu/shift_result[25] ) );
BUF_X1 \malu/Shift/_1532_ ( .A(\malu/Shift/_0739_ ), .Z(\malu/shift_result[26] ) );
BUF_X1 \malu/Shift/_1533_ ( .A(\malu/Shift/_0740_ ), .Z(\malu/shift_result[27] ) );
BUF_X1 \malu/Shift/_1534_ ( .A(\malu/Shift/_0741_ ), .Z(\malu/shift_result[28] ) );
BUF_X1 \malu/Shift/_1535_ ( .A(\malu/Shift/_0742_ ), .Z(\malu/shift_result[29] ) );
BUF_X1 \malu/Shift/_1536_ ( .A(\malu/Shift/_0744_ ), .Z(\malu/shift_result[30] ) );
BUF_X1 \malu/Shift/_1537_ ( .A(\malu/Shift/_0745_ ), .Z(\malu/shift_result[31] ) );
NAND2_X4 \marbiter/_0710_ ( .A1(\marbiter/_0702_ ), .A2(\marbiter/_0214_ ), .ZN(\marbiter/_0228_ ) );
INV_X8 \marbiter/_0711_ ( .A(\marbiter/_0571_ ), .ZN(\marbiter/_0229_ ) );
NAND3_X1 \marbiter/_0712_ ( .A1(\marbiter/_0228_ ), .A2(\marbiter/_0229_ ), .A3(\marbiter/_0674_ ), .ZN(\marbiter/_0230_ ) );
AND2_X4 \marbiter/_0713_ ( .A1(\marbiter/_0703_ ), .A2(\marbiter/_0215_ ), .ZN(\marbiter/_0231_ ) );
NOR2_X1 \marbiter/_0714_ ( .A1(\marbiter/_0230_ ), .A2(\marbiter/_0231_ ), .ZN(\marbiter/_0232_ ) );
AND2_X2 \marbiter/_0715_ ( .A1(\marbiter/_0671_ ), .A2(\marbiter/_0676_ ), .ZN(\marbiter/_0672_ ) );
AND2_X4 \marbiter/_0716_ ( .A1(\marbiter/_0671_ ), .A2(\marbiter/_0675_ ), .ZN(\marbiter/_0673_ ) );
OR4_X2 \marbiter/_0717_ ( .A1(\marbiter/_0571_ ), .A2(\marbiter/_0232_ ), .A3(\marbiter/_0672_ ), .A4(\marbiter/_0673_ ), .ZN(\marbiter/_0009_ ) );
NAND3_X1 \marbiter/_0718_ ( .A1(\marbiter/_0229_ ), .A2(\marbiter/_0112_ ), .A3(\marbiter/_0559_ ), .ZN(\marbiter/_0233_ ) );
OR2_X1 \marbiter/_0719_ ( .A1(\marbiter/_0571_ ), .A2(\marbiter/_0572_ ), .ZN(\marbiter/_0234_ ) );
INV_X1 \marbiter/_0720_ ( .A(\marbiter/_0561_ ), .ZN(\marbiter/_0235_ ) );
OAI21_X1 \marbiter/_0721_ ( .A(\marbiter/_0233_ ), .B1(\marbiter/_0234_ ), .B2(\marbiter/_0235_ ), .ZN(\marbiter/_0008_ ) );
NAND4_X1 \marbiter/_0722_ ( .A1(\marbiter/_0231_ ), .A2(\marbiter/_0229_ ), .A3(\marbiter/_0674_ ), .A4(\marbiter/_0228_ ), .ZN(\marbiter/_0236_ ) );
INV_X1 \marbiter/_0723_ ( .A(\marbiter/_0675_ ), .ZN(\marbiter/_0237_ ) );
OR2_X1 \marbiter/_0724_ ( .A1(\marbiter/_0571_ ), .A2(\marbiter/_0671_ ), .ZN(\marbiter/_0238_ ) );
OAI21_X1 \marbiter/_0725_ ( .A(\marbiter/_0236_ ), .B1(\marbiter/_0237_ ), .B2(\marbiter/_0238_ ), .ZN(\marbiter/_0010_ ) );
NAND4_X1 \marbiter/_0726_ ( .A1(\marbiter/_0229_ ), .A2(\marbiter/_0702_ ), .A3(\marbiter/_0214_ ), .A4(\marbiter/_0674_ ), .ZN(\marbiter/_0239_ ) );
INV_X1 \marbiter/_0727_ ( .A(\marbiter/_0676_ ), .ZN(\marbiter/_0240_ ) );
OAI21_X1 \marbiter/_0728_ ( .A(\marbiter/_0239_ ), .B1(\marbiter/_0238_ ), .B2(\marbiter/_0240_ ), .ZN(\marbiter/_0011_ ) );
NOR3_X1 \marbiter/_0729_ ( .A1(\marbiter/_0571_ ), .A2(\marbiter/_0112_ ), .A3(\marbiter/_0113_ ), .ZN(\marbiter/_0241_ ) );
AND2_X1 \marbiter/_0730_ ( .A1(\marbiter/_0241_ ), .A2(\marbiter/_0559_ ), .ZN(\marbiter/_0242_ ) );
AND2_X2 \marbiter/_0731_ ( .A1(\marbiter/_0572_ ), .A2(\marbiter/_0560_ ), .ZN(\marbiter/_0574_ ) );
AND2_X4 \marbiter/_0732_ ( .A1(\marbiter/_0572_ ), .A2(\marbiter/_0561_ ), .ZN(\marbiter/_0573_ ) );
OR4_X2 \marbiter/_0733_ ( .A1(\marbiter/_0571_ ), .A2(\marbiter/_0242_ ), .A3(\marbiter/_0574_ ), .A4(\marbiter/_0573_ ), .ZN(\marbiter/_0006_ ) );
INV_X1 \marbiter/_0734_ ( .A(\marbiter/_0112_ ), .ZN(\marbiter/_0243_ ) );
NAND4_X1 \marbiter/_0735_ ( .A1(\marbiter/_0229_ ), .A2(\marbiter/_0243_ ), .A3(\marbiter/_0559_ ), .A4(\marbiter/_0113_ ), .ZN(\marbiter/_0244_ ) );
INV_X1 \marbiter/_0736_ ( .A(\marbiter/_0560_ ), .ZN(\marbiter/_0245_ ) );
OAI21_X1 \marbiter/_0737_ ( .A(\marbiter/_0244_ ), .B1(\marbiter/_0245_ ), .B2(\marbiter/_0234_ ), .ZN(\marbiter/_0007_ ) );
AND2_X1 \marbiter/_0738_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0569_ ), .ZN(\marbiter/_0565_ ) );
AND2_X1 \marbiter/_0739_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0570_ ), .ZN(\marbiter/_0566_ ) );
AND2_X1 \marbiter/_0740_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0527_ ), .ZN(\marbiter/_0463_ ) );
AND2_X1 \marbiter/_0741_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0538_ ), .ZN(\marbiter/_0474_ ) );
AND2_X1 \marbiter/_0742_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0549_ ), .ZN(\marbiter/_0485_ ) );
AND2_X1 \marbiter/_0743_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0552_ ), .ZN(\marbiter/_0488_ ) );
AND2_X1 \marbiter/_0744_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0553_ ), .ZN(\marbiter/_0489_ ) );
AND2_X1 \marbiter/_0745_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0554_ ), .ZN(\marbiter/_0490_ ) );
AND2_X1 \marbiter/_0746_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0555_ ), .ZN(\marbiter/_0491_ ) );
AND2_X1 \marbiter/_0747_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0556_ ), .ZN(\marbiter/_0492_ ) );
AND2_X1 \marbiter/_0748_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0557_ ), .ZN(\marbiter/_0493_ ) );
AND2_X1 \marbiter/_0749_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0558_ ), .ZN(\marbiter/_0494_ ) );
AND2_X1 \marbiter/_0750_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0528_ ), .ZN(\marbiter/_0464_ ) );
AND2_X1 \marbiter/_0751_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0529_ ), .ZN(\marbiter/_0465_ ) );
AND2_X1 \marbiter/_0752_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0530_ ), .ZN(\marbiter/_0466_ ) );
AND2_X1 \marbiter/_0753_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0531_ ), .ZN(\marbiter/_0467_ ) );
AND2_X1 \marbiter/_0754_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0532_ ), .ZN(\marbiter/_0468_ ) );
AND2_X1 \marbiter/_0755_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0533_ ), .ZN(\marbiter/_0469_ ) );
AND2_X1 \marbiter/_0756_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0534_ ), .ZN(\marbiter/_0470_ ) );
AND2_X1 \marbiter/_0757_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0535_ ), .ZN(\marbiter/_0471_ ) );
AND2_X1 \marbiter/_0758_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0536_ ), .ZN(\marbiter/_0472_ ) );
AND2_X1 \marbiter/_0759_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0537_ ), .ZN(\marbiter/_0473_ ) );
AND2_X1 \marbiter/_0760_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0539_ ), .ZN(\marbiter/_0475_ ) );
AND2_X1 \marbiter/_0761_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0540_ ), .ZN(\marbiter/_0476_ ) );
AND2_X1 \marbiter/_0762_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0541_ ), .ZN(\marbiter/_0477_ ) );
AND2_X1 \marbiter/_0763_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0542_ ), .ZN(\marbiter/_0478_ ) );
AND2_X1 \marbiter/_0764_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0543_ ), .ZN(\marbiter/_0479_ ) );
AND2_X1 \marbiter/_0765_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0544_ ), .ZN(\marbiter/_0480_ ) );
AND2_X1 \marbiter/_0766_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0545_ ), .ZN(\marbiter/_0481_ ) );
AND2_X1 \marbiter/_0767_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0546_ ), .ZN(\marbiter/_0482_ ) );
AND2_X1 \marbiter/_0768_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0547_ ), .ZN(\marbiter/_0483_ ) );
AND2_X1 \marbiter/_0769_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0548_ ), .ZN(\marbiter/_0484_ ) );
AND2_X1 \marbiter/_0770_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0550_ ), .ZN(\marbiter/_0486_ ) );
AND2_X1 \marbiter/_0771_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0551_ ), .ZN(\marbiter/_0487_ ) );
AND2_X1 \marbiter/_0772_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0569_ ), .ZN(\marbiter/_0567_ ) );
AND2_X1 \marbiter/_0773_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0570_ ), .ZN(\marbiter/_0568_ ) );
AND2_X1 \marbiter/_0774_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0527_ ), .ZN(\marbiter/_0495_ ) );
AND2_X1 \marbiter/_0775_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0538_ ), .ZN(\marbiter/_0506_ ) );
AND2_X1 \marbiter/_0776_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0549_ ), .ZN(\marbiter/_0517_ ) );
AND2_X1 \marbiter/_0777_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0552_ ), .ZN(\marbiter/_0520_ ) );
AND2_X1 \marbiter/_0778_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0553_ ), .ZN(\marbiter/_0521_ ) );
AND2_X1 \marbiter/_0779_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0554_ ), .ZN(\marbiter/_0522_ ) );
AND2_X1 \marbiter/_0780_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0555_ ), .ZN(\marbiter/_0523_ ) );
AND2_X1 \marbiter/_0781_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0556_ ), .ZN(\marbiter/_0524_ ) );
AND2_X1 \marbiter/_0782_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0557_ ), .ZN(\marbiter/_0525_ ) );
AND2_X1 \marbiter/_0783_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0558_ ), .ZN(\marbiter/_0526_ ) );
AND2_X1 \marbiter/_0784_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0528_ ), .ZN(\marbiter/_0496_ ) );
AND2_X1 \marbiter/_0785_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0529_ ), .ZN(\marbiter/_0497_ ) );
AND2_X1 \marbiter/_0786_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0530_ ), .ZN(\marbiter/_0498_ ) );
AND2_X1 \marbiter/_0787_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0531_ ), .ZN(\marbiter/_0499_ ) );
AND2_X1 \marbiter/_0788_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0532_ ), .ZN(\marbiter/_0500_ ) );
AND2_X1 \marbiter/_0789_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0533_ ), .ZN(\marbiter/_0501_ ) );
AND2_X1 \marbiter/_0790_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0534_ ), .ZN(\marbiter/_0502_ ) );
AND2_X1 \marbiter/_0791_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0535_ ), .ZN(\marbiter/_0503_ ) );
AND2_X1 \marbiter/_0792_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0536_ ), .ZN(\marbiter/_0504_ ) );
AND2_X1 \marbiter/_0793_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0537_ ), .ZN(\marbiter/_0505_ ) );
AND2_X1 \marbiter/_0794_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0539_ ), .ZN(\marbiter/_0507_ ) );
AND2_X1 \marbiter/_0795_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0540_ ), .ZN(\marbiter/_0508_ ) );
AND2_X1 \marbiter/_0796_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0541_ ), .ZN(\marbiter/_0509_ ) );
AND2_X1 \marbiter/_0797_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0542_ ), .ZN(\marbiter/_0510_ ) );
AND2_X1 \marbiter/_0798_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0543_ ), .ZN(\marbiter/_0511_ ) );
AND2_X1 \marbiter/_0799_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0544_ ), .ZN(\marbiter/_0512_ ) );
AND2_X1 \marbiter/_0800_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0545_ ), .ZN(\marbiter/_0513_ ) );
AND2_X1 \marbiter/_0801_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0546_ ), .ZN(\marbiter/_0514_ ) );
AND2_X1 \marbiter/_0802_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0547_ ), .ZN(\marbiter/_0515_ ) );
AND2_X1 \marbiter/_0803_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0548_ ), .ZN(\marbiter/_0516_ ) );
AND2_X1 \marbiter/_0804_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0550_ ), .ZN(\marbiter/_0518_ ) );
AND2_X1 \marbiter/_0805_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0551_ ), .ZN(\marbiter/_0519_ ) );
AND2_X1 \marbiter/_0806_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0223_ ), .ZN(\marbiter/_0219_ ) );
AND2_X1 \marbiter/_0807_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0224_ ), .ZN(\marbiter/_0220_ ) );
AND2_X1 \marbiter/_0808_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0223_ ), .ZN(\marbiter/_0221_ ) );
AND2_X1 \marbiter/_0809_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0224_ ), .ZN(\marbiter/_0222_ ) );
NAND2_X1 \marbiter/_0810_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0685_ ), .ZN(\marbiter/_0246_ ) );
NAND2_X1 \marbiter/_0811_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0677_ ), .ZN(\marbiter/_0247_ ) );
NAND2_X1 \marbiter/_0812_ ( .A1(\marbiter/_0246_ ), .A2(\marbiter/_0247_ ), .ZN(\marbiter/_0693_ ) );
NAND2_X1 \marbiter/_0813_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0686_ ), .ZN(\marbiter/_0248_ ) );
NAND2_X1 \marbiter/_0814_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0678_ ), .ZN(\marbiter/_0249_ ) );
NAND2_X1 \marbiter/_0815_ ( .A1(\marbiter/_0248_ ), .A2(\marbiter/_0249_ ), .ZN(\marbiter/_0694_ ) );
NAND2_X1 \marbiter/_0816_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0687_ ), .ZN(\marbiter/_0250_ ) );
NAND2_X1 \marbiter/_0817_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0679_ ), .ZN(\marbiter/_0251_ ) );
NAND2_X1 \marbiter/_0818_ ( .A1(\marbiter/_0250_ ), .A2(\marbiter/_0251_ ), .ZN(\marbiter/_0695_ ) );
NAND2_X1 \marbiter/_0819_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0688_ ), .ZN(\marbiter/_0252_ ) );
NAND2_X1 \marbiter/_0820_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0680_ ), .ZN(\marbiter/_0253_ ) );
NAND2_X1 \marbiter/_0821_ ( .A1(\marbiter/_0252_ ), .A2(\marbiter/_0253_ ), .ZN(\marbiter/_0696_ ) );
NAND2_X1 \marbiter/_0822_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0689_ ), .ZN(\marbiter/_0254_ ) );
NAND2_X1 \marbiter/_0823_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0681_ ), .ZN(\marbiter/_0255_ ) );
NAND2_X1 \marbiter/_0824_ ( .A1(\marbiter/_0254_ ), .A2(\marbiter/_0255_ ), .ZN(\marbiter/_0697_ ) );
NAND2_X1 \marbiter/_0825_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0690_ ), .ZN(\marbiter/_0256_ ) );
NAND2_X1 \marbiter/_0826_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0682_ ), .ZN(\marbiter/_0257_ ) );
NAND2_X1 \marbiter/_0827_ ( .A1(\marbiter/_0256_ ), .A2(\marbiter/_0257_ ), .ZN(\marbiter/_0698_ ) );
NAND2_X1 \marbiter/_0828_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0691_ ), .ZN(\marbiter/_0258_ ) );
NAND2_X1 \marbiter/_0829_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0683_ ), .ZN(\marbiter/_0259_ ) );
NAND2_X1 \marbiter/_0830_ ( .A1(\marbiter/_0258_ ), .A2(\marbiter/_0259_ ), .ZN(\marbiter/_0699_ ) );
NAND2_X1 \marbiter/_0831_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0692_ ), .ZN(\marbiter/_0260_ ) );
NAND2_X1 \marbiter/_0832_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0684_ ), .ZN(\marbiter/_0261_ ) );
NAND2_X1 \marbiter/_0833_ ( .A1(\marbiter/_0260_ ), .A2(\marbiter/_0261_ ), .ZN(\marbiter/_0700_ ) );
NAND2_X1 \marbiter/_0834_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0607_ ), .ZN(\marbiter/_0262_ ) );
NAND2_X1 \marbiter/_0835_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0575_ ), .ZN(\marbiter/_0263_ ) );
NAND2_X1 \marbiter/_0836_ ( .A1(\marbiter/_0262_ ), .A2(\marbiter/_0263_ ), .ZN(\marbiter/_0639_ ) );
NAND2_X1 \marbiter/_0837_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0618_ ), .ZN(\marbiter/_0264_ ) );
NAND2_X1 \marbiter/_0838_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0586_ ), .ZN(\marbiter/_0265_ ) );
NAND2_X1 \marbiter/_0839_ ( .A1(\marbiter/_0264_ ), .A2(\marbiter/_0265_ ), .ZN(\marbiter/_0650_ ) );
NAND2_X1 \marbiter/_0840_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0629_ ), .ZN(\marbiter/_0266_ ) );
NAND2_X1 \marbiter/_0841_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0597_ ), .ZN(\marbiter/_0267_ ) );
NAND2_X1 \marbiter/_0842_ ( .A1(\marbiter/_0266_ ), .A2(\marbiter/_0267_ ), .ZN(\marbiter/_0661_ ) );
NAND2_X1 \marbiter/_0843_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0632_ ), .ZN(\marbiter/_0268_ ) );
NAND2_X1 \marbiter/_0844_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0600_ ), .ZN(\marbiter/_0269_ ) );
NAND2_X1 \marbiter/_0845_ ( .A1(\marbiter/_0268_ ), .A2(\marbiter/_0269_ ), .ZN(\marbiter/_0664_ ) );
NAND2_X1 \marbiter/_0846_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0633_ ), .ZN(\marbiter/_0270_ ) );
NAND2_X1 \marbiter/_0847_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0601_ ), .ZN(\marbiter/_0271_ ) );
NAND2_X1 \marbiter/_0848_ ( .A1(\marbiter/_0270_ ), .A2(\marbiter/_0271_ ), .ZN(\marbiter/_0665_ ) );
NAND2_X1 \marbiter/_0849_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0634_ ), .ZN(\marbiter/_0272_ ) );
NAND2_X1 \marbiter/_0850_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0602_ ), .ZN(\marbiter/_0273_ ) );
NAND2_X1 \marbiter/_0851_ ( .A1(\marbiter/_0272_ ), .A2(\marbiter/_0273_ ), .ZN(\marbiter/_0666_ ) );
NAND2_X1 \marbiter/_0852_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0635_ ), .ZN(\marbiter/_0274_ ) );
NAND2_X1 \marbiter/_0853_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0603_ ), .ZN(\marbiter/_0275_ ) );
NAND2_X1 \marbiter/_0854_ ( .A1(\marbiter/_0274_ ), .A2(\marbiter/_0275_ ), .ZN(\marbiter/_0667_ ) );
NAND2_X1 \marbiter/_0855_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0636_ ), .ZN(\marbiter/_0276_ ) );
NAND2_X1 \marbiter/_0856_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0604_ ), .ZN(\marbiter/_0277_ ) );
NAND2_X1 \marbiter/_0857_ ( .A1(\marbiter/_0276_ ), .A2(\marbiter/_0277_ ), .ZN(\marbiter/_0668_ ) );
NAND2_X1 \marbiter/_0858_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0637_ ), .ZN(\marbiter/_0278_ ) );
NAND2_X1 \marbiter/_0859_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0605_ ), .ZN(\marbiter/_0279_ ) );
NAND2_X1 \marbiter/_0860_ ( .A1(\marbiter/_0278_ ), .A2(\marbiter/_0279_ ), .ZN(\marbiter/_0669_ ) );
NAND2_X1 \marbiter/_0861_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0638_ ), .ZN(\marbiter/_0280_ ) );
NAND2_X1 \marbiter/_0862_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0606_ ), .ZN(\marbiter/_0281_ ) );
NAND2_X1 \marbiter/_0863_ ( .A1(\marbiter/_0280_ ), .A2(\marbiter/_0281_ ), .ZN(\marbiter/_0670_ ) );
NAND2_X1 \marbiter/_0864_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0608_ ), .ZN(\marbiter/_0282_ ) );
NAND2_X1 \marbiter/_0865_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0576_ ), .ZN(\marbiter/_0283_ ) );
NAND2_X1 \marbiter/_0866_ ( .A1(\marbiter/_0282_ ), .A2(\marbiter/_0283_ ), .ZN(\marbiter/_0640_ ) );
NAND2_X1 \marbiter/_0867_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0609_ ), .ZN(\marbiter/_0284_ ) );
NAND2_X1 \marbiter/_0868_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0577_ ), .ZN(\marbiter/_0285_ ) );
NAND2_X1 \marbiter/_0869_ ( .A1(\marbiter/_0284_ ), .A2(\marbiter/_0285_ ), .ZN(\marbiter/_0641_ ) );
NAND2_X1 \marbiter/_0870_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0610_ ), .ZN(\marbiter/_0286_ ) );
NAND2_X1 \marbiter/_0871_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0578_ ), .ZN(\marbiter/_0287_ ) );
NAND2_X1 \marbiter/_0872_ ( .A1(\marbiter/_0286_ ), .A2(\marbiter/_0287_ ), .ZN(\marbiter/_0642_ ) );
NAND2_X1 \marbiter/_0873_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0611_ ), .ZN(\marbiter/_0288_ ) );
NAND2_X1 \marbiter/_0874_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0579_ ), .ZN(\marbiter/_0289_ ) );
NAND2_X1 \marbiter/_0875_ ( .A1(\marbiter/_0288_ ), .A2(\marbiter/_0289_ ), .ZN(\marbiter/_0643_ ) );
NAND2_X1 \marbiter/_0876_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0612_ ), .ZN(\marbiter/_0290_ ) );
NAND2_X1 \marbiter/_0877_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0580_ ), .ZN(\marbiter/_0291_ ) );
NAND2_X1 \marbiter/_0878_ ( .A1(\marbiter/_0290_ ), .A2(\marbiter/_0291_ ), .ZN(\marbiter/_0644_ ) );
NAND2_X1 \marbiter/_0879_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0613_ ), .ZN(\marbiter/_0292_ ) );
NAND2_X1 \marbiter/_0880_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0581_ ), .ZN(\marbiter/_0293_ ) );
NAND2_X1 \marbiter/_0881_ ( .A1(\marbiter/_0292_ ), .A2(\marbiter/_0293_ ), .ZN(\marbiter/_0645_ ) );
NAND2_X1 \marbiter/_0882_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0614_ ), .ZN(\marbiter/_0294_ ) );
NAND2_X1 \marbiter/_0883_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0582_ ), .ZN(\marbiter/_0295_ ) );
NAND2_X1 \marbiter/_0884_ ( .A1(\marbiter/_0294_ ), .A2(\marbiter/_0295_ ), .ZN(\marbiter/_0646_ ) );
NAND2_X1 \marbiter/_0885_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0615_ ), .ZN(\marbiter/_0296_ ) );
NAND2_X1 \marbiter/_0886_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0583_ ), .ZN(\marbiter/_0297_ ) );
NAND2_X1 \marbiter/_0887_ ( .A1(\marbiter/_0296_ ), .A2(\marbiter/_0297_ ), .ZN(\marbiter/_0647_ ) );
NAND2_X1 \marbiter/_0888_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0616_ ), .ZN(\marbiter/_0298_ ) );
NAND2_X1 \marbiter/_0889_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0584_ ), .ZN(\marbiter/_0299_ ) );
NAND2_X1 \marbiter/_0890_ ( .A1(\marbiter/_0298_ ), .A2(\marbiter/_0299_ ), .ZN(\marbiter/_0648_ ) );
NAND2_X1 \marbiter/_0891_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0617_ ), .ZN(\marbiter/_0300_ ) );
NAND2_X1 \marbiter/_0892_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0585_ ), .ZN(\marbiter/_0301_ ) );
NAND2_X1 \marbiter/_0893_ ( .A1(\marbiter/_0300_ ), .A2(\marbiter/_0301_ ), .ZN(\marbiter/_0649_ ) );
NAND2_X1 \marbiter/_0894_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0619_ ), .ZN(\marbiter/_0302_ ) );
NAND2_X1 \marbiter/_0895_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0587_ ), .ZN(\marbiter/_0303_ ) );
NAND2_X1 \marbiter/_0896_ ( .A1(\marbiter/_0302_ ), .A2(\marbiter/_0303_ ), .ZN(\marbiter/_0651_ ) );
NAND2_X1 \marbiter/_0897_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0620_ ), .ZN(\marbiter/_0304_ ) );
NAND2_X1 \marbiter/_0898_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0588_ ), .ZN(\marbiter/_0305_ ) );
NAND2_X1 \marbiter/_0899_ ( .A1(\marbiter/_0304_ ), .A2(\marbiter/_0305_ ), .ZN(\marbiter/_0652_ ) );
NAND2_X1 \marbiter/_0900_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0621_ ), .ZN(\marbiter/_0306_ ) );
NAND2_X1 \marbiter/_0901_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0589_ ), .ZN(\marbiter/_0307_ ) );
NAND2_X1 \marbiter/_0902_ ( .A1(\marbiter/_0306_ ), .A2(\marbiter/_0307_ ), .ZN(\marbiter/_0653_ ) );
NAND2_X1 \marbiter/_0903_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0622_ ), .ZN(\marbiter/_0308_ ) );
NAND2_X1 \marbiter/_0904_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0590_ ), .ZN(\marbiter/_0309_ ) );
NAND2_X1 \marbiter/_0905_ ( .A1(\marbiter/_0308_ ), .A2(\marbiter/_0309_ ), .ZN(\marbiter/_0654_ ) );
NAND2_X1 \marbiter/_0906_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0623_ ), .ZN(\marbiter/_0310_ ) );
NAND2_X1 \marbiter/_0907_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0591_ ), .ZN(\marbiter/_0311_ ) );
NAND2_X1 \marbiter/_0908_ ( .A1(\marbiter/_0310_ ), .A2(\marbiter/_0311_ ), .ZN(\marbiter/_0655_ ) );
NAND2_X1 \marbiter/_0909_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0624_ ), .ZN(\marbiter/_0312_ ) );
NAND2_X1 \marbiter/_0910_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0592_ ), .ZN(\marbiter/_0313_ ) );
NAND2_X1 \marbiter/_0911_ ( .A1(\marbiter/_0312_ ), .A2(\marbiter/_0313_ ), .ZN(\marbiter/_0656_ ) );
NAND2_X1 \marbiter/_0912_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0625_ ), .ZN(\marbiter/_0314_ ) );
NAND2_X1 \marbiter/_0913_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0593_ ), .ZN(\marbiter/_0315_ ) );
NAND2_X1 \marbiter/_0914_ ( .A1(\marbiter/_0314_ ), .A2(\marbiter/_0315_ ), .ZN(\marbiter/_0657_ ) );
NAND2_X1 \marbiter/_0915_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0626_ ), .ZN(\marbiter/_0316_ ) );
NAND2_X1 \marbiter/_0916_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0594_ ), .ZN(\marbiter/_0317_ ) );
NAND2_X1 \marbiter/_0917_ ( .A1(\marbiter/_0316_ ), .A2(\marbiter/_0317_ ), .ZN(\marbiter/_0658_ ) );
NAND2_X1 \marbiter/_0918_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0627_ ), .ZN(\marbiter/_0318_ ) );
NAND2_X1 \marbiter/_0919_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0595_ ), .ZN(\marbiter/_0319_ ) );
NAND2_X1 \marbiter/_0920_ ( .A1(\marbiter/_0318_ ), .A2(\marbiter/_0319_ ), .ZN(\marbiter/_0659_ ) );
NAND2_X1 \marbiter/_0921_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0628_ ), .ZN(\marbiter/_0320_ ) );
NAND2_X1 \marbiter/_0922_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0596_ ), .ZN(\marbiter/_0321_ ) );
NAND2_X1 \marbiter/_0923_ ( .A1(\marbiter/_0320_ ), .A2(\marbiter/_0321_ ), .ZN(\marbiter/_0660_ ) );
NAND2_X1 \marbiter/_0924_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0630_ ), .ZN(\marbiter/_0322_ ) );
NAND2_X1 \marbiter/_0925_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0598_ ), .ZN(\marbiter/_0323_ ) );
NAND2_X1 \marbiter/_0926_ ( .A1(\marbiter/_0322_ ), .A2(\marbiter/_0323_ ), .ZN(\marbiter/_0662_ ) );
NAND2_X1 \marbiter/_0927_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0631_ ), .ZN(\marbiter/_0324_ ) );
NAND2_X1 \marbiter/_0928_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0599_ ), .ZN(\marbiter/_0325_ ) );
NAND2_X1 \marbiter/_0929_ ( .A1(\marbiter/_0324_ ), .A2(\marbiter/_0325_ ), .ZN(\marbiter/_0663_ ) );
NAND2_X1 \marbiter/_0930_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0146_ ), .ZN(\marbiter/_0326_ ) );
NAND2_X1 \marbiter/_0931_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0114_ ), .ZN(\marbiter/_0327_ ) );
NAND2_X1 \marbiter/_0932_ ( .A1(\marbiter/_0326_ ), .A2(\marbiter/_0327_ ), .ZN(\marbiter/_0178_ ) );
NAND2_X1 \marbiter/_0933_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0157_ ), .ZN(\marbiter/_0328_ ) );
NAND2_X1 \marbiter/_0934_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0125_ ), .ZN(\marbiter/_0329_ ) );
NAND2_X1 \marbiter/_0935_ ( .A1(\marbiter/_0328_ ), .A2(\marbiter/_0329_ ), .ZN(\marbiter/_0189_ ) );
NAND2_X1 \marbiter/_0936_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0168_ ), .ZN(\marbiter/_0330_ ) );
NAND2_X1 \marbiter/_0937_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0136_ ), .ZN(\marbiter/_0331_ ) );
NAND2_X1 \marbiter/_0938_ ( .A1(\marbiter/_0330_ ), .A2(\marbiter/_0331_ ), .ZN(\marbiter/_0200_ ) );
NAND2_X1 \marbiter/_0939_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0171_ ), .ZN(\marbiter/_0332_ ) );
NAND2_X1 \marbiter/_0940_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0139_ ), .ZN(\marbiter/_0333_ ) );
NAND2_X1 \marbiter/_0941_ ( .A1(\marbiter/_0332_ ), .A2(\marbiter/_0333_ ), .ZN(\marbiter/_0203_ ) );
NAND2_X1 \marbiter/_0942_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0172_ ), .ZN(\marbiter/_0334_ ) );
NAND2_X1 \marbiter/_0943_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0140_ ), .ZN(\marbiter/_0335_ ) );
NAND2_X1 \marbiter/_0944_ ( .A1(\marbiter/_0334_ ), .A2(\marbiter/_0335_ ), .ZN(\marbiter/_0204_ ) );
NAND2_X1 \marbiter/_0945_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0173_ ), .ZN(\marbiter/_0336_ ) );
NAND2_X1 \marbiter/_0946_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0141_ ), .ZN(\marbiter/_0337_ ) );
NAND2_X1 \marbiter/_0947_ ( .A1(\marbiter/_0336_ ), .A2(\marbiter/_0337_ ), .ZN(\marbiter/_0205_ ) );
NAND2_X1 \marbiter/_0948_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0174_ ), .ZN(\marbiter/_0338_ ) );
NAND2_X1 \marbiter/_0949_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0142_ ), .ZN(\marbiter/_0339_ ) );
NAND2_X1 \marbiter/_0950_ ( .A1(\marbiter/_0338_ ), .A2(\marbiter/_0339_ ), .ZN(\marbiter/_0206_ ) );
NAND2_X1 \marbiter/_0951_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0175_ ), .ZN(\marbiter/_0340_ ) );
NAND2_X1 \marbiter/_0952_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0143_ ), .ZN(\marbiter/_0341_ ) );
NAND2_X1 \marbiter/_0953_ ( .A1(\marbiter/_0340_ ), .A2(\marbiter/_0341_ ), .ZN(\marbiter/_0207_ ) );
NAND2_X1 \marbiter/_0954_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0176_ ), .ZN(\marbiter/_0342_ ) );
NAND2_X1 \marbiter/_0955_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0144_ ), .ZN(\marbiter/_0343_ ) );
NAND2_X1 \marbiter/_0956_ ( .A1(\marbiter/_0342_ ), .A2(\marbiter/_0343_ ), .ZN(\marbiter/_0208_ ) );
NAND2_X1 \marbiter/_0957_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0177_ ), .ZN(\marbiter/_0344_ ) );
NAND2_X1 \marbiter/_0958_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0145_ ), .ZN(\marbiter/_0345_ ) );
NAND2_X1 \marbiter/_0959_ ( .A1(\marbiter/_0344_ ), .A2(\marbiter/_0345_ ), .ZN(\marbiter/_0209_ ) );
NAND2_X1 \marbiter/_0960_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0147_ ), .ZN(\marbiter/_0346_ ) );
NAND2_X1 \marbiter/_0961_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0115_ ), .ZN(\marbiter/_0347_ ) );
NAND2_X1 \marbiter/_0962_ ( .A1(\marbiter/_0346_ ), .A2(\marbiter/_0347_ ), .ZN(\marbiter/_0179_ ) );
NAND2_X1 \marbiter/_0963_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0148_ ), .ZN(\marbiter/_0348_ ) );
NAND2_X1 \marbiter/_0964_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0116_ ), .ZN(\marbiter/_0349_ ) );
NAND2_X1 \marbiter/_0965_ ( .A1(\marbiter/_0348_ ), .A2(\marbiter/_0349_ ), .ZN(\marbiter/_0180_ ) );
NAND2_X1 \marbiter/_0966_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0149_ ), .ZN(\marbiter/_0350_ ) );
NAND2_X1 \marbiter/_0967_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0117_ ), .ZN(\marbiter/_0351_ ) );
NAND2_X1 \marbiter/_0968_ ( .A1(\marbiter/_0350_ ), .A2(\marbiter/_0351_ ), .ZN(\marbiter/_0181_ ) );
NAND2_X1 \marbiter/_0969_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0150_ ), .ZN(\marbiter/_0352_ ) );
NAND2_X1 \marbiter/_0970_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0118_ ), .ZN(\marbiter/_0353_ ) );
NAND2_X1 \marbiter/_0971_ ( .A1(\marbiter/_0352_ ), .A2(\marbiter/_0353_ ), .ZN(\marbiter/_0182_ ) );
NAND2_X1 \marbiter/_0972_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0151_ ), .ZN(\marbiter/_0354_ ) );
NAND2_X1 \marbiter/_0973_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0119_ ), .ZN(\marbiter/_0355_ ) );
NAND2_X1 \marbiter/_0974_ ( .A1(\marbiter/_0354_ ), .A2(\marbiter/_0355_ ), .ZN(\marbiter/_0183_ ) );
NAND2_X1 \marbiter/_0975_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0152_ ), .ZN(\marbiter/_0356_ ) );
NAND2_X1 \marbiter/_0976_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0120_ ), .ZN(\marbiter/_0357_ ) );
NAND2_X1 \marbiter/_0977_ ( .A1(\marbiter/_0356_ ), .A2(\marbiter/_0357_ ), .ZN(\marbiter/_0184_ ) );
NAND2_X1 \marbiter/_0978_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0153_ ), .ZN(\marbiter/_0358_ ) );
NAND2_X1 \marbiter/_0979_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0121_ ), .ZN(\marbiter/_0359_ ) );
NAND2_X1 \marbiter/_0980_ ( .A1(\marbiter/_0358_ ), .A2(\marbiter/_0359_ ), .ZN(\marbiter/_0185_ ) );
NAND2_X1 \marbiter/_0981_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0154_ ), .ZN(\marbiter/_0360_ ) );
NAND2_X1 \marbiter/_0982_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0122_ ), .ZN(\marbiter/_0361_ ) );
NAND2_X1 \marbiter/_0983_ ( .A1(\marbiter/_0360_ ), .A2(\marbiter/_0361_ ), .ZN(\marbiter/_0186_ ) );
NAND2_X1 \marbiter/_0984_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0155_ ), .ZN(\marbiter/_0362_ ) );
NAND2_X1 \marbiter/_0985_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0123_ ), .ZN(\marbiter/_0363_ ) );
NAND2_X1 \marbiter/_0986_ ( .A1(\marbiter/_0362_ ), .A2(\marbiter/_0363_ ), .ZN(\marbiter/_0187_ ) );
NAND2_X1 \marbiter/_0987_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0156_ ), .ZN(\marbiter/_0364_ ) );
NAND2_X1 \marbiter/_0988_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0124_ ), .ZN(\marbiter/_0365_ ) );
NAND2_X1 \marbiter/_0989_ ( .A1(\marbiter/_0364_ ), .A2(\marbiter/_0365_ ), .ZN(\marbiter/_0188_ ) );
NAND2_X1 \marbiter/_0990_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0158_ ), .ZN(\marbiter/_0366_ ) );
NAND2_X1 \marbiter/_0991_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0126_ ), .ZN(\marbiter/_0367_ ) );
NAND2_X1 \marbiter/_0992_ ( .A1(\marbiter/_0366_ ), .A2(\marbiter/_0367_ ), .ZN(\marbiter/_0190_ ) );
NAND2_X1 \marbiter/_0993_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0159_ ), .ZN(\marbiter/_0368_ ) );
NAND2_X1 \marbiter/_0994_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0127_ ), .ZN(\marbiter/_0369_ ) );
NAND2_X1 \marbiter/_0995_ ( .A1(\marbiter/_0368_ ), .A2(\marbiter/_0369_ ), .ZN(\marbiter/_0191_ ) );
NAND2_X1 \marbiter/_0996_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0160_ ), .ZN(\marbiter/_0370_ ) );
NAND2_X1 \marbiter/_0997_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0128_ ), .ZN(\marbiter/_0371_ ) );
NAND2_X1 \marbiter/_0998_ ( .A1(\marbiter/_0370_ ), .A2(\marbiter/_0371_ ), .ZN(\marbiter/_0192_ ) );
NAND2_X1 \marbiter/_0999_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0161_ ), .ZN(\marbiter/_0372_ ) );
NAND2_X1 \marbiter/_1000_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0129_ ), .ZN(\marbiter/_0373_ ) );
NAND2_X1 \marbiter/_1001_ ( .A1(\marbiter/_0372_ ), .A2(\marbiter/_0373_ ), .ZN(\marbiter/_0193_ ) );
NAND2_X1 \marbiter/_1002_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0162_ ), .ZN(\marbiter/_0374_ ) );
NAND2_X1 \marbiter/_1003_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0130_ ), .ZN(\marbiter/_0375_ ) );
NAND2_X1 \marbiter/_1004_ ( .A1(\marbiter/_0374_ ), .A2(\marbiter/_0375_ ), .ZN(\marbiter/_0194_ ) );
NAND2_X1 \marbiter/_1005_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0163_ ), .ZN(\marbiter/_0376_ ) );
NAND2_X1 \marbiter/_1006_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0131_ ), .ZN(\marbiter/_0377_ ) );
NAND2_X1 \marbiter/_1007_ ( .A1(\marbiter/_0376_ ), .A2(\marbiter/_0377_ ), .ZN(\marbiter/_0195_ ) );
NAND2_X1 \marbiter/_1008_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0164_ ), .ZN(\marbiter/_0378_ ) );
NAND2_X1 \marbiter/_1009_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0132_ ), .ZN(\marbiter/_0379_ ) );
NAND2_X1 \marbiter/_1010_ ( .A1(\marbiter/_0378_ ), .A2(\marbiter/_0379_ ), .ZN(\marbiter/_0196_ ) );
NAND2_X1 \marbiter/_1011_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0165_ ), .ZN(\marbiter/_0380_ ) );
NAND2_X1 \marbiter/_1012_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0133_ ), .ZN(\marbiter/_0381_ ) );
NAND2_X1 \marbiter/_1013_ ( .A1(\marbiter/_0380_ ), .A2(\marbiter/_0381_ ), .ZN(\marbiter/_0197_ ) );
NAND2_X1 \marbiter/_1014_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0166_ ), .ZN(\marbiter/_0382_ ) );
NAND2_X1 \marbiter/_1015_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0134_ ), .ZN(\marbiter/_0383_ ) );
NAND2_X1 \marbiter/_1016_ ( .A1(\marbiter/_0382_ ), .A2(\marbiter/_0383_ ), .ZN(\marbiter/_0198_ ) );
NAND2_X1 \marbiter/_1017_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0167_ ), .ZN(\marbiter/_0384_ ) );
NAND2_X1 \marbiter/_1018_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0135_ ), .ZN(\marbiter/_0385_ ) );
NAND2_X1 \marbiter/_1019_ ( .A1(\marbiter/_0384_ ), .A2(\marbiter/_0385_ ), .ZN(\marbiter/_0199_ ) );
NAND2_X1 \marbiter/_1020_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0169_ ), .ZN(\marbiter/_0386_ ) );
NAND2_X1 \marbiter/_1021_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0137_ ), .ZN(\marbiter/_0387_ ) );
NAND2_X1 \marbiter/_1022_ ( .A1(\marbiter/_0386_ ), .A2(\marbiter/_0387_ ), .ZN(\marbiter/_0201_ ) );
NAND2_X1 \marbiter/_1023_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0170_ ), .ZN(\marbiter/_0388_ ) );
NAND2_X1 \marbiter/_1024_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0138_ ), .ZN(\marbiter/_0389_ ) );
NAND2_X1 \marbiter/_1025_ ( .A1(\marbiter/_0388_ ), .A2(\marbiter/_0389_ ), .ZN(\marbiter/_0202_ ) );
NAND2_X1 \marbiter/_1026_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0218_ ), .ZN(\marbiter/_0390_ ) );
NAND2_X1 \marbiter/_1027_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0217_ ), .ZN(\marbiter/_0391_ ) );
NAND2_X1 \marbiter/_1028_ ( .A1(\marbiter/_0390_ ), .A2(\marbiter/_0391_ ), .ZN(\marbiter/_0216_ ) );
NAND2_X1 \marbiter/_1029_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0703_ ), .ZN(\marbiter/_0392_ ) );
NAND2_X1 \marbiter/_1030_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0702_ ), .ZN(\marbiter/_0393_ ) );
NAND2_X1 \marbiter/_1031_ ( .A1(\marbiter/_0392_ ), .A2(\marbiter/_0393_ ), .ZN(\marbiter/_0701_ ) );
NAND2_X1 \marbiter/_1032_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0215_ ), .ZN(\marbiter/_0394_ ) );
NAND2_X1 \marbiter/_1033_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0214_ ), .ZN(\marbiter/_0395_ ) );
NAND2_X1 \marbiter/_1034_ ( .A1(\marbiter/_0394_ ), .A2(\marbiter/_0395_ ), .ZN(\marbiter/_0213_ ) );
NAND2_X1 \marbiter/_1035_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0044_ ), .ZN(\marbiter/_0396_ ) );
NAND2_X1 \marbiter/_1036_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0012_ ), .ZN(\marbiter/_0397_ ) );
NAND2_X1 \marbiter/_1037_ ( .A1(\marbiter/_0396_ ), .A2(\marbiter/_0397_ ), .ZN(\marbiter/_0076_ ) );
NAND2_X1 \marbiter/_1038_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0055_ ), .ZN(\marbiter/_0398_ ) );
NAND2_X1 \marbiter/_1039_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0023_ ), .ZN(\marbiter/_0399_ ) );
NAND2_X1 \marbiter/_1040_ ( .A1(\marbiter/_0398_ ), .A2(\marbiter/_0399_ ), .ZN(\marbiter/_0087_ ) );
NAND2_X1 \marbiter/_1041_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0066_ ), .ZN(\marbiter/_0400_ ) );
NAND2_X1 \marbiter/_1042_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0034_ ), .ZN(\marbiter/_0401_ ) );
NAND2_X1 \marbiter/_1043_ ( .A1(\marbiter/_0400_ ), .A2(\marbiter/_0401_ ), .ZN(\marbiter/_0098_ ) );
NAND2_X1 \marbiter/_1044_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0069_ ), .ZN(\marbiter/_0402_ ) );
NAND2_X1 \marbiter/_1045_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0037_ ), .ZN(\marbiter/_0403_ ) );
NAND2_X1 \marbiter/_1046_ ( .A1(\marbiter/_0402_ ), .A2(\marbiter/_0403_ ), .ZN(\marbiter/_0101_ ) );
NAND2_X1 \marbiter/_1047_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0070_ ), .ZN(\marbiter/_0404_ ) );
NAND2_X1 \marbiter/_1048_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0038_ ), .ZN(\marbiter/_0405_ ) );
NAND2_X1 \marbiter/_1049_ ( .A1(\marbiter/_0404_ ), .A2(\marbiter/_0405_ ), .ZN(\marbiter/_0102_ ) );
NAND2_X1 \marbiter/_1050_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0071_ ), .ZN(\marbiter/_0406_ ) );
NAND2_X1 \marbiter/_1051_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0039_ ), .ZN(\marbiter/_0407_ ) );
NAND2_X1 \marbiter/_1052_ ( .A1(\marbiter/_0406_ ), .A2(\marbiter/_0407_ ), .ZN(\marbiter/_0103_ ) );
NAND2_X1 \marbiter/_1053_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0072_ ), .ZN(\marbiter/_0408_ ) );
NAND2_X1 \marbiter/_1054_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0040_ ), .ZN(\marbiter/_0409_ ) );
NAND2_X1 \marbiter/_1055_ ( .A1(\marbiter/_0408_ ), .A2(\marbiter/_0409_ ), .ZN(\marbiter/_0104_ ) );
NAND2_X1 \marbiter/_1056_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0073_ ), .ZN(\marbiter/_0410_ ) );
NAND2_X1 \marbiter/_1057_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0041_ ), .ZN(\marbiter/_0411_ ) );
NAND2_X1 \marbiter/_1058_ ( .A1(\marbiter/_0410_ ), .A2(\marbiter/_0411_ ), .ZN(\marbiter/_0105_ ) );
NAND2_X1 \marbiter/_1059_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0074_ ), .ZN(\marbiter/_0412_ ) );
NAND2_X1 \marbiter/_1060_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0042_ ), .ZN(\marbiter/_0413_ ) );
NAND2_X1 \marbiter/_1061_ ( .A1(\marbiter/_0412_ ), .A2(\marbiter/_0413_ ), .ZN(\marbiter/_0106_ ) );
NAND2_X1 \marbiter/_1062_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0075_ ), .ZN(\marbiter/_0414_ ) );
NAND2_X1 \marbiter/_1063_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0043_ ), .ZN(\marbiter/_0415_ ) );
NAND2_X1 \marbiter/_1064_ ( .A1(\marbiter/_0414_ ), .A2(\marbiter/_0415_ ), .ZN(\marbiter/_0107_ ) );
NAND2_X1 \marbiter/_1065_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0045_ ), .ZN(\marbiter/_0416_ ) );
NAND2_X1 \marbiter/_1066_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0013_ ), .ZN(\marbiter/_0417_ ) );
NAND2_X1 \marbiter/_1067_ ( .A1(\marbiter/_0416_ ), .A2(\marbiter/_0417_ ), .ZN(\marbiter/_0077_ ) );
NAND2_X1 \marbiter/_1068_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0046_ ), .ZN(\marbiter/_0418_ ) );
NAND2_X1 \marbiter/_1069_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0014_ ), .ZN(\marbiter/_0419_ ) );
NAND2_X1 \marbiter/_1070_ ( .A1(\marbiter/_0418_ ), .A2(\marbiter/_0419_ ), .ZN(\marbiter/_0078_ ) );
NAND2_X1 \marbiter/_1071_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0047_ ), .ZN(\marbiter/_0420_ ) );
NAND2_X1 \marbiter/_1072_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0015_ ), .ZN(\marbiter/_0421_ ) );
NAND2_X1 \marbiter/_1073_ ( .A1(\marbiter/_0420_ ), .A2(\marbiter/_0421_ ), .ZN(\marbiter/_0079_ ) );
NAND2_X1 \marbiter/_1074_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0048_ ), .ZN(\marbiter/_0422_ ) );
NAND2_X1 \marbiter/_1075_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0016_ ), .ZN(\marbiter/_0423_ ) );
NAND2_X1 \marbiter/_1076_ ( .A1(\marbiter/_0422_ ), .A2(\marbiter/_0423_ ), .ZN(\marbiter/_0080_ ) );
NAND2_X1 \marbiter/_1077_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0049_ ), .ZN(\marbiter/_0424_ ) );
NAND2_X1 \marbiter/_1078_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0017_ ), .ZN(\marbiter/_0425_ ) );
NAND2_X1 \marbiter/_1079_ ( .A1(\marbiter/_0424_ ), .A2(\marbiter/_0425_ ), .ZN(\marbiter/_0081_ ) );
NAND2_X1 \marbiter/_1080_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0050_ ), .ZN(\marbiter/_0426_ ) );
NAND2_X1 \marbiter/_1081_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0018_ ), .ZN(\marbiter/_0427_ ) );
NAND2_X1 \marbiter/_1082_ ( .A1(\marbiter/_0426_ ), .A2(\marbiter/_0427_ ), .ZN(\marbiter/_0082_ ) );
NAND2_X1 \marbiter/_1083_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0051_ ), .ZN(\marbiter/_0428_ ) );
NAND2_X1 \marbiter/_1084_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0019_ ), .ZN(\marbiter/_0429_ ) );
NAND2_X1 \marbiter/_1085_ ( .A1(\marbiter/_0428_ ), .A2(\marbiter/_0429_ ), .ZN(\marbiter/_0083_ ) );
NAND2_X1 \marbiter/_1086_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0052_ ), .ZN(\marbiter/_0430_ ) );
NAND2_X1 \marbiter/_1087_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0020_ ), .ZN(\marbiter/_0431_ ) );
NAND2_X1 \marbiter/_1088_ ( .A1(\marbiter/_0430_ ), .A2(\marbiter/_0431_ ), .ZN(\marbiter/_0084_ ) );
NAND2_X1 \marbiter/_1089_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0053_ ), .ZN(\marbiter/_0432_ ) );
NAND2_X1 \marbiter/_1090_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0021_ ), .ZN(\marbiter/_0433_ ) );
NAND2_X1 \marbiter/_1091_ ( .A1(\marbiter/_0432_ ), .A2(\marbiter/_0433_ ), .ZN(\marbiter/_0085_ ) );
NAND2_X1 \marbiter/_1092_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0054_ ), .ZN(\marbiter/_0434_ ) );
NAND2_X1 \marbiter/_1093_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0022_ ), .ZN(\marbiter/_0435_ ) );
NAND2_X1 \marbiter/_1094_ ( .A1(\marbiter/_0434_ ), .A2(\marbiter/_0435_ ), .ZN(\marbiter/_0086_ ) );
NAND2_X1 \marbiter/_1095_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0056_ ), .ZN(\marbiter/_0436_ ) );
NAND2_X1 \marbiter/_1096_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0024_ ), .ZN(\marbiter/_0437_ ) );
NAND2_X1 \marbiter/_1097_ ( .A1(\marbiter/_0436_ ), .A2(\marbiter/_0437_ ), .ZN(\marbiter/_0088_ ) );
NAND2_X1 \marbiter/_1098_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0057_ ), .ZN(\marbiter/_0438_ ) );
NAND2_X1 \marbiter/_1099_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0025_ ), .ZN(\marbiter/_0439_ ) );
NAND2_X1 \marbiter/_1100_ ( .A1(\marbiter/_0438_ ), .A2(\marbiter/_0439_ ), .ZN(\marbiter/_0089_ ) );
NAND2_X1 \marbiter/_1101_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0058_ ), .ZN(\marbiter/_0440_ ) );
NAND2_X1 \marbiter/_1102_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0026_ ), .ZN(\marbiter/_0441_ ) );
NAND2_X1 \marbiter/_1103_ ( .A1(\marbiter/_0440_ ), .A2(\marbiter/_0441_ ), .ZN(\marbiter/_0090_ ) );
NAND2_X1 \marbiter/_1104_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0059_ ), .ZN(\marbiter/_0442_ ) );
NAND2_X1 \marbiter/_1105_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0027_ ), .ZN(\marbiter/_0443_ ) );
NAND2_X1 \marbiter/_1106_ ( .A1(\marbiter/_0442_ ), .A2(\marbiter/_0443_ ), .ZN(\marbiter/_0091_ ) );
NAND2_X1 \marbiter/_1107_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0060_ ), .ZN(\marbiter/_0444_ ) );
NAND2_X1 \marbiter/_1108_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0028_ ), .ZN(\marbiter/_0445_ ) );
NAND2_X1 \marbiter/_1109_ ( .A1(\marbiter/_0444_ ), .A2(\marbiter/_0445_ ), .ZN(\marbiter/_0092_ ) );
NAND2_X1 \marbiter/_1110_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0061_ ), .ZN(\marbiter/_0446_ ) );
NAND2_X1 \marbiter/_1111_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0029_ ), .ZN(\marbiter/_0447_ ) );
NAND2_X1 \marbiter/_1112_ ( .A1(\marbiter/_0446_ ), .A2(\marbiter/_0447_ ), .ZN(\marbiter/_0093_ ) );
NAND2_X1 \marbiter/_1113_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0062_ ), .ZN(\marbiter/_0448_ ) );
NAND2_X1 \marbiter/_1114_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0030_ ), .ZN(\marbiter/_0449_ ) );
NAND2_X1 \marbiter/_1115_ ( .A1(\marbiter/_0448_ ), .A2(\marbiter/_0449_ ), .ZN(\marbiter/_0094_ ) );
NAND2_X1 \marbiter/_1116_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0063_ ), .ZN(\marbiter/_0450_ ) );
NAND2_X1 \marbiter/_1117_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0031_ ), .ZN(\marbiter/_0451_ ) );
NAND2_X1 \marbiter/_1118_ ( .A1(\marbiter/_0450_ ), .A2(\marbiter/_0451_ ), .ZN(\marbiter/_0095_ ) );
NAND2_X1 \marbiter/_1119_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0064_ ), .ZN(\marbiter/_0452_ ) );
NAND2_X1 \marbiter/_1120_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0032_ ), .ZN(\marbiter/_0453_ ) );
NAND2_X1 \marbiter/_1121_ ( .A1(\marbiter/_0452_ ), .A2(\marbiter/_0453_ ), .ZN(\marbiter/_0096_ ) );
NAND2_X1 \marbiter/_1122_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0065_ ), .ZN(\marbiter/_0454_ ) );
NAND2_X1 \marbiter/_1123_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0033_ ), .ZN(\marbiter/_0455_ ) );
NAND2_X1 \marbiter/_1124_ ( .A1(\marbiter/_0454_ ), .A2(\marbiter/_0455_ ), .ZN(\marbiter/_0097_ ) );
NAND2_X1 \marbiter/_1125_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0067_ ), .ZN(\marbiter/_0456_ ) );
NAND2_X1 \marbiter/_1126_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0035_ ), .ZN(\marbiter/_0457_ ) );
NAND2_X1 \marbiter/_1127_ ( .A1(\marbiter/_0456_ ), .A2(\marbiter/_0457_ ), .ZN(\marbiter/_0099_ ) );
NAND2_X1 \marbiter/_1128_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0068_ ), .ZN(\marbiter/_0458_ ) );
NAND2_X1 \marbiter/_1129_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0036_ ), .ZN(\marbiter/_0459_ ) );
NAND2_X1 \marbiter/_1130_ ( .A1(\marbiter/_0458_ ), .A2(\marbiter/_0459_ ), .ZN(\marbiter/_0100_ ) );
NAND2_X1 \marbiter/_1131_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0564_ ), .ZN(\marbiter/_0460_ ) );
NAND2_X1 \marbiter/_1132_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0563_ ), .ZN(\marbiter/_0461_ ) );
NAND2_X1 \marbiter/_1133_ ( .A1(\marbiter/_0460_ ), .A2(\marbiter/_0461_ ), .ZN(\marbiter/_0562_ ) );
NAND2_X1 \marbiter/_1134_ ( .A1(\marbiter/_0113_ ), .A2(\marbiter/_0560_ ), .ZN(\marbiter/_0462_ ) );
OAI21_X1 \marbiter/_1135_ ( .A(\marbiter/_0462_ ), .B1(\marbiter/_0243_ ), .B2(\marbiter/_0235_ ), .ZN(\marbiter/_0111_ ) );
AND2_X1 \marbiter/_1136_ ( .A1(\marbiter/_0561_ ), .A2(\marbiter/_0108_ ), .ZN(\marbiter/_0109_ ) );
AND2_X1 \marbiter/_1137_ ( .A1(\marbiter/_0560_ ), .A2(\marbiter/_0108_ ), .ZN(\marbiter/_0110_ ) );
AND2_X1 \marbiter/_1138_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0210_ ), .ZN(\marbiter/_0211_ ) );
AND2_X1 \marbiter/_1139_ ( .A1(\marbiter/_0676_ ), .A2(\marbiter/_0225_ ), .ZN(\marbiter/_0226_ ) );
AND2_X1 \marbiter/_1140_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0210_ ), .ZN(\marbiter/_0212_ ) );
AND2_X1 \marbiter/_1141_ ( .A1(\marbiter/_0675_ ), .A2(\marbiter/_0225_ ), .ZN(\marbiter/_0227_ ) );
DFF_X1 \marbiter/_1142_ ( .CK(clk ), .D(\marbiter/_0003_ ), .Q(\marbiter/write_state[0] ), .QN(\marbiter/_0705_ ) );
DFF_X1 \marbiter/_1143_ ( .CK(clk ), .D(\marbiter/_0004_ ), .Q(\marbiter/write_state[1] ), .QN(\marbiter/_0706_ ) );
DFF_X1 \marbiter/_1144_ ( .CK(clk ), .D(\marbiter/_0005_ ), .Q(\marbiter/write_state[2] ), .QN(\marbiter/_0707_ ) );
DFF_X1 \marbiter/_1145_ ( .CK(clk ), .D(\marbiter/_0000_ ), .Q(\marbiter/read_state[0] ), .QN(\marbiter/_0708_ ) );
DFF_X1 \marbiter/_1146_ ( .CK(clk ), .D(\marbiter/_0001_ ), .Q(\marbiter/read_state[1] ), .QN(\marbiter/_0709_ ) );
DFF_X1 \marbiter/_1147_ ( .CK(clk ), .D(\marbiter/_0002_ ), .Q(\marbiter/read_state[2] ), .QN(\marbiter/_0704_ ) );
BUF_X1 \marbiter/_1148_ ( .A(rst ), .Z(\marbiter/_0571_ ) );
BUF_X1 \marbiter/_1149_ ( .A(wready ), .Z(\marbiter/_0671_ ) );
BUF_X1 \marbiter/_1150_ ( .A(\marbiter/write_state[2] ), .Z(\marbiter/_0676_ ) );
BUF_X1 \marbiter/_1151_ ( .A(\marbiter/write_state[1] ), .Z(\marbiter/_0675_ ) );
BUF_X1 \marbiter/_1152_ ( .A(_351_ ), .Z(\marbiter/_0702_ ) );
BUF_X1 \marbiter/_1153_ ( .A(_351_ ), .Z(\marbiter/_0214_ ) );
BUF_X1 \marbiter/_1154_ ( .A(lsu_wvalid ), .Z(\marbiter/_0703_ ) );
BUF_X1 \marbiter/_1155_ ( .A(lsu_awvalid ), .Z(\marbiter/_0215_ ) );
BUF_X1 \marbiter/_1156_ ( .A(\marbiter/write_state[0] ), .Z(\marbiter/_0674_ ) );
BUF_X1 \marbiter/_1157_ ( .A(\marbiter/_0009_ ), .Z(\marbiter/_0003_ ) );
BUF_X1 \marbiter/_1158_ ( .A(ifu_arvalid ), .Z(\marbiter/_0112_ ) );
BUF_X1 \marbiter/_1159_ ( .A(\marbiter/read_state[0] ), .Z(\marbiter/_0559_ ) );
BUF_X1 \marbiter/_1160_ ( .A(rvalid ), .Z(\marbiter/_0572_ ) );
BUF_X1 \marbiter/_1161_ ( .A(\marbiter/read_state[2] ), .Z(\marbiter/_0561_ ) );
BUF_X1 \marbiter/_1162_ ( .A(\marbiter/_0008_ ), .Z(\marbiter/_0002_ ) );
BUF_X1 \marbiter/_1163_ ( .A(\marbiter/_0010_ ), .Z(\marbiter/_0004_ ) );
BUF_X1 \marbiter/_1164_ ( .A(\marbiter/_0011_ ), .Z(\marbiter/_0005_ ) );
BUF_X1 \marbiter/_1165_ ( .A(lsu_arvalid ), .Z(\marbiter/_0113_ ) );
BUF_X1 \marbiter/_1166_ ( .A(\marbiter/read_state[1] ), .Z(\marbiter/_0560_ ) );
BUF_X1 \marbiter/_1167_ ( .A(\marbiter/_0006_ ), .Z(\marbiter/_0000_ ) );
BUF_X1 \marbiter/_1168_ ( .A(\marbiter/_0007_ ), .Z(\marbiter/_0001_ ) );
BUF_X1 \marbiter/_1169_ ( .A(\rresp[0] ), .Z(\marbiter/_0569_ ) );
BUF_X1 \marbiter/_1170_ ( .A(\marbiter/_0565_ ), .Z(\ifu_rresp[0] ) );
BUF_X1 \marbiter/_1171_ ( .A(\rresp[1] ), .Z(\marbiter/_0570_ ) );
BUF_X1 \marbiter/_1172_ ( .A(\marbiter/_0566_ ), .Z(\ifu_rresp[1] ) );
BUF_X1 \marbiter/_1173_ ( .A(\rdata[0] ), .Z(\marbiter/_0527_ ) );
BUF_X1 \marbiter/_1174_ ( .A(\marbiter/_0463_ ), .Z(\ifu_rdata[0] ) );
BUF_X1 \marbiter/_1175_ ( .A(\rdata[1] ), .Z(\marbiter/_0538_ ) );
BUF_X1 \marbiter/_1176_ ( .A(\marbiter/_0474_ ), .Z(\ifu_rdata[1] ) );
BUF_X1 \marbiter/_1177_ ( .A(\rdata[2] ), .Z(\marbiter/_0549_ ) );
BUF_X1 \marbiter/_1178_ ( .A(\marbiter/_0485_ ), .Z(\ifu_rdata[2] ) );
BUF_X1 \marbiter/_1179_ ( .A(\rdata[3] ), .Z(\marbiter/_0552_ ) );
BUF_X1 \marbiter/_1180_ ( .A(\marbiter/_0488_ ), .Z(\ifu_rdata[3] ) );
BUF_X1 \marbiter/_1181_ ( .A(\rdata[4] ), .Z(\marbiter/_0553_ ) );
BUF_X1 \marbiter/_1182_ ( .A(\marbiter/_0489_ ), .Z(\ifu_rdata[4] ) );
BUF_X1 \marbiter/_1183_ ( .A(\rdata[5] ), .Z(\marbiter/_0554_ ) );
BUF_X1 \marbiter/_1184_ ( .A(\marbiter/_0490_ ), .Z(\ifu_rdata[5] ) );
BUF_X1 \marbiter/_1185_ ( .A(\rdata[6] ), .Z(\marbiter/_0555_ ) );
BUF_X1 \marbiter/_1186_ ( .A(\marbiter/_0491_ ), .Z(\ifu_rdata[6] ) );
BUF_X1 \marbiter/_1187_ ( .A(\rdata[7] ), .Z(\marbiter/_0556_ ) );
BUF_X1 \marbiter/_1188_ ( .A(\marbiter/_0492_ ), .Z(\ifu_rdata[7] ) );
BUF_X1 \marbiter/_1189_ ( .A(\rdata[8] ), .Z(\marbiter/_0557_ ) );
BUF_X1 \marbiter/_1190_ ( .A(\marbiter/_0493_ ), .Z(\ifu_rdata[8] ) );
BUF_X1 \marbiter/_1191_ ( .A(\rdata[9] ), .Z(\marbiter/_0558_ ) );
BUF_X1 \marbiter/_1192_ ( .A(\marbiter/_0494_ ), .Z(\ifu_rdata[9] ) );
BUF_X1 \marbiter/_1193_ ( .A(\rdata[10] ), .Z(\marbiter/_0528_ ) );
BUF_X1 \marbiter/_1194_ ( .A(\marbiter/_0464_ ), .Z(\ifu_rdata[10] ) );
BUF_X1 \marbiter/_1195_ ( .A(\rdata[11] ), .Z(\marbiter/_0529_ ) );
BUF_X1 \marbiter/_1196_ ( .A(\marbiter/_0465_ ), .Z(\ifu_rdata[11] ) );
BUF_X1 \marbiter/_1197_ ( .A(\rdata[12] ), .Z(\marbiter/_0530_ ) );
BUF_X1 \marbiter/_1198_ ( .A(\marbiter/_0466_ ), .Z(\ifu_rdata[12] ) );
BUF_X1 \marbiter/_1199_ ( .A(\rdata[13] ), .Z(\marbiter/_0531_ ) );
BUF_X1 \marbiter/_1200_ ( .A(\marbiter/_0467_ ), .Z(\ifu_rdata[13] ) );
BUF_X1 \marbiter/_1201_ ( .A(\rdata[14] ), .Z(\marbiter/_0532_ ) );
BUF_X1 \marbiter/_1202_ ( .A(\marbiter/_0468_ ), .Z(\ifu_rdata[14] ) );
BUF_X1 \marbiter/_1203_ ( .A(\rdata[15] ), .Z(\marbiter/_0533_ ) );
BUF_X1 \marbiter/_1204_ ( .A(\marbiter/_0469_ ), .Z(\ifu_rdata[15] ) );
BUF_X1 \marbiter/_1205_ ( .A(\rdata[16] ), .Z(\marbiter/_0534_ ) );
BUF_X1 \marbiter/_1206_ ( .A(\marbiter/_0470_ ), .Z(\ifu_rdata[16] ) );
BUF_X1 \marbiter/_1207_ ( .A(\rdata[17] ), .Z(\marbiter/_0535_ ) );
BUF_X1 \marbiter/_1208_ ( .A(\marbiter/_0471_ ), .Z(\ifu_rdata[17] ) );
BUF_X1 \marbiter/_1209_ ( .A(\rdata[18] ), .Z(\marbiter/_0536_ ) );
BUF_X1 \marbiter/_1210_ ( .A(\marbiter/_0472_ ), .Z(\ifu_rdata[18] ) );
BUF_X1 \marbiter/_1211_ ( .A(\rdata[19] ), .Z(\marbiter/_0537_ ) );
BUF_X1 \marbiter/_1212_ ( .A(\marbiter/_0473_ ), .Z(\ifu_rdata[19] ) );
BUF_X1 \marbiter/_1213_ ( .A(\rdata[20] ), .Z(\marbiter/_0539_ ) );
BUF_X1 \marbiter/_1214_ ( .A(\marbiter/_0475_ ), .Z(\ifu_rdata[20] ) );
BUF_X1 \marbiter/_1215_ ( .A(\rdata[21] ), .Z(\marbiter/_0540_ ) );
BUF_X1 \marbiter/_1216_ ( .A(\marbiter/_0476_ ), .Z(\ifu_rdata[21] ) );
BUF_X1 \marbiter/_1217_ ( .A(\rdata[22] ), .Z(\marbiter/_0541_ ) );
BUF_X1 \marbiter/_1218_ ( .A(\marbiter/_0477_ ), .Z(\ifu_rdata[22] ) );
BUF_X1 \marbiter/_1219_ ( .A(\rdata[23] ), .Z(\marbiter/_0542_ ) );
BUF_X1 \marbiter/_1220_ ( .A(\marbiter/_0478_ ), .Z(\ifu_rdata[23] ) );
BUF_X1 \marbiter/_1221_ ( .A(\rdata[24] ), .Z(\marbiter/_0543_ ) );
BUF_X1 \marbiter/_1222_ ( .A(\marbiter/_0479_ ), .Z(\ifu_rdata[24] ) );
BUF_X1 \marbiter/_1223_ ( .A(\rdata[25] ), .Z(\marbiter/_0544_ ) );
BUF_X1 \marbiter/_1224_ ( .A(\marbiter/_0480_ ), .Z(\ifu_rdata[25] ) );
BUF_X1 \marbiter/_1225_ ( .A(\rdata[26] ), .Z(\marbiter/_0545_ ) );
BUF_X1 \marbiter/_1226_ ( .A(\marbiter/_0481_ ), .Z(\ifu_rdata[26] ) );
BUF_X1 \marbiter/_1227_ ( .A(\rdata[27] ), .Z(\marbiter/_0546_ ) );
BUF_X1 \marbiter/_1228_ ( .A(\marbiter/_0482_ ), .Z(\ifu_rdata[27] ) );
BUF_X1 \marbiter/_1229_ ( .A(\rdata[28] ), .Z(\marbiter/_0547_ ) );
BUF_X1 \marbiter/_1230_ ( .A(\marbiter/_0483_ ), .Z(\ifu_rdata[28] ) );
BUF_X1 \marbiter/_1231_ ( .A(\rdata[29] ), .Z(\marbiter/_0548_ ) );
BUF_X1 \marbiter/_1232_ ( .A(\marbiter/_0484_ ), .Z(\ifu_rdata[29] ) );
BUF_X1 \marbiter/_1233_ ( .A(\rdata[30] ), .Z(\marbiter/_0550_ ) );
BUF_X1 \marbiter/_1234_ ( .A(\marbiter/_0486_ ), .Z(\ifu_rdata[30] ) );
BUF_X1 \marbiter/_1235_ ( .A(\rdata[31] ), .Z(\marbiter/_0551_ ) );
BUF_X1 \marbiter/_1236_ ( .A(\marbiter/_0487_ ), .Z(\ifu_rdata[31] ) );
BUF_X1 \marbiter/_1237_ ( .A(\marbiter/_0567_ ), .Z(\lsu_rresp[0] ) );
BUF_X1 \marbiter/_1238_ ( .A(\marbiter/_0568_ ), .Z(\lsu_rresp[1] ) );
BUF_X1 \marbiter/_1239_ ( .A(\marbiter/_0495_ ), .Z(\lsu_rdata[0] ) );
BUF_X1 \marbiter/_1240_ ( .A(\marbiter/_0506_ ), .Z(\lsu_rdata[1] ) );
BUF_X1 \marbiter/_1241_ ( .A(\marbiter/_0517_ ), .Z(\lsu_rdata[2] ) );
BUF_X1 \marbiter/_1242_ ( .A(\marbiter/_0520_ ), .Z(\lsu_rdata[3] ) );
BUF_X1 \marbiter/_1243_ ( .A(\marbiter/_0521_ ), .Z(\lsu_rdata[4] ) );
BUF_X1 \marbiter/_1244_ ( .A(\marbiter/_0522_ ), .Z(\lsu_rdata[5] ) );
BUF_X1 \marbiter/_1245_ ( .A(\marbiter/_0523_ ), .Z(\lsu_rdata[6] ) );
BUF_X1 \marbiter/_1246_ ( .A(\marbiter/_0524_ ), .Z(\lsu_rdata[7] ) );
BUF_X1 \marbiter/_1247_ ( .A(\marbiter/_0525_ ), .Z(\lsu_rdata[8] ) );
BUF_X1 \marbiter/_1248_ ( .A(\marbiter/_0526_ ), .Z(\lsu_rdata[9] ) );
BUF_X1 \marbiter/_1249_ ( .A(\marbiter/_0496_ ), .Z(\lsu_rdata[10] ) );
BUF_X1 \marbiter/_1250_ ( .A(\marbiter/_0497_ ), .Z(\lsu_rdata[11] ) );
BUF_X1 \marbiter/_1251_ ( .A(\marbiter/_0498_ ), .Z(\lsu_rdata[12] ) );
BUF_X1 \marbiter/_1252_ ( .A(\marbiter/_0499_ ), .Z(\lsu_rdata[13] ) );
BUF_X1 \marbiter/_1253_ ( .A(\marbiter/_0500_ ), .Z(\lsu_rdata[14] ) );
BUF_X1 \marbiter/_1254_ ( .A(\marbiter/_0501_ ), .Z(\lsu_rdata[15] ) );
BUF_X1 \marbiter/_1255_ ( .A(\marbiter/_0502_ ), .Z(\lsu_rdata[16] ) );
BUF_X1 \marbiter/_1256_ ( .A(\marbiter/_0503_ ), .Z(\lsu_rdata[17] ) );
BUF_X1 \marbiter/_1257_ ( .A(\marbiter/_0504_ ), .Z(\lsu_rdata[18] ) );
BUF_X1 \marbiter/_1258_ ( .A(\marbiter/_0505_ ), .Z(\lsu_rdata[19] ) );
BUF_X1 \marbiter/_1259_ ( .A(\marbiter/_0507_ ), .Z(\lsu_rdata[20] ) );
BUF_X1 \marbiter/_1260_ ( .A(\marbiter/_0508_ ), .Z(\lsu_rdata[21] ) );
BUF_X1 \marbiter/_1261_ ( .A(\marbiter/_0509_ ), .Z(\lsu_rdata[22] ) );
BUF_X1 \marbiter/_1262_ ( .A(\marbiter/_0510_ ), .Z(\lsu_rdata[23] ) );
BUF_X1 \marbiter/_1263_ ( .A(\marbiter/_0511_ ), .Z(\lsu_rdata[24] ) );
BUF_X1 \marbiter/_1264_ ( .A(\marbiter/_0512_ ), .Z(\lsu_rdata[25] ) );
BUF_X1 \marbiter/_1265_ ( .A(\marbiter/_0513_ ), .Z(\lsu_rdata[26] ) );
BUF_X1 \marbiter/_1266_ ( .A(\marbiter/_0514_ ), .Z(\lsu_rdata[27] ) );
BUF_X1 \marbiter/_1267_ ( .A(\marbiter/_0515_ ), .Z(\lsu_rdata[28] ) );
BUF_X1 \marbiter/_1268_ ( .A(\marbiter/_0516_ ), .Z(\lsu_rdata[29] ) );
BUF_X1 \marbiter/_1269_ ( .A(\marbiter/_0518_ ), .Z(\lsu_rdata[30] ) );
BUF_X1 \marbiter/_1270_ ( .A(\marbiter/_0519_ ), .Z(\lsu_rdata[31] ) );
BUF_X1 \marbiter/_1271_ ( .A(\bresp[0] ), .Z(\marbiter/_0223_ ) );
BUF_X1 \marbiter/_1272_ ( .A(\marbiter/_0219_ ), .Z(\ifu_bresp[0] ) );
BUF_X1 \marbiter/_1273_ ( .A(\bresp[1] ), .Z(\marbiter/_0224_ ) );
BUF_X1 \marbiter/_1274_ ( .A(\marbiter/_0220_ ), .Z(\ifu_bresp[1] ) );
BUF_X1 \marbiter/_1275_ ( .A(\marbiter/_0221_ ), .Z(\lsu_bresp[0] ) );
BUF_X1 \marbiter/_1276_ ( .A(\marbiter/_0222_ ), .Z(\lsu_bresp[1] ) );
BUF_X1 \marbiter/_1277_ ( .A(\lsu_wstrb[0] ), .Z(\marbiter/_0685_ ) );
BUF_X1 \marbiter/_1278_ ( .A(_351_ ), .Z(\marbiter/_0677_ ) );
BUF_X1 \marbiter/_1279_ ( .A(\marbiter/_0693_ ), .Z(\wstrb[0] ) );
BUF_X1 \marbiter/_1280_ ( .A(\lsu_wstrb[1] ), .Z(\marbiter/_0686_ ) );
BUF_X1 \marbiter/_1281_ ( .A(_351_ ), .Z(\marbiter/_0678_ ) );
BUF_X1 \marbiter/_1282_ ( .A(\marbiter/_0694_ ), .Z(\wstrb[1] ) );
BUF_X1 \marbiter/_1283_ ( .A(\lsu_wstrb[2] ), .Z(\marbiter/_0687_ ) );
BUF_X1 \marbiter/_1284_ ( .A(_351_ ), .Z(\marbiter/_0679_ ) );
BUF_X1 \marbiter/_1285_ ( .A(\marbiter/_0695_ ), .Z(\wstrb[2] ) );
BUF_X1 \marbiter/_1286_ ( .A(\lsu_wstrb[3] ), .Z(\marbiter/_0688_ ) );
BUF_X1 \marbiter/_1287_ ( .A(_351_ ), .Z(\marbiter/_0680_ ) );
BUF_X1 \marbiter/_1288_ ( .A(\marbiter/_0696_ ), .Z(\wstrb[3] ) );
BUF_X1 \marbiter/_1289_ ( .A(\lsu_wstrb[4] ), .Z(\marbiter/_0689_ ) );
BUF_X1 \marbiter/_1290_ ( .A(_351_ ), .Z(\marbiter/_0681_ ) );
BUF_X1 \marbiter/_1291_ ( .A(\marbiter/_0697_ ), .Z(\wstrb[4] ) );
BUF_X1 \marbiter/_1292_ ( .A(\lsu_wstrb[5] ), .Z(\marbiter/_0690_ ) );
BUF_X1 \marbiter/_1293_ ( .A(_351_ ), .Z(\marbiter/_0682_ ) );
BUF_X1 \marbiter/_1294_ ( .A(\marbiter/_0698_ ), .Z(\wstrb[5] ) );
BUF_X1 \marbiter/_1295_ ( .A(\lsu_wstrb[6] ), .Z(\marbiter/_0691_ ) );
BUF_X1 \marbiter/_1296_ ( .A(_351_ ), .Z(\marbiter/_0683_ ) );
BUF_X1 \marbiter/_1297_ ( .A(\marbiter/_0699_ ), .Z(\wstrb[6] ) );
BUF_X1 \marbiter/_1298_ ( .A(\lsu_wstrb[7] ), .Z(\marbiter/_0692_ ) );
BUF_X1 \marbiter/_1299_ ( .A(_351_ ), .Z(\marbiter/_0684_ ) );
BUF_X1 \marbiter/_1300_ ( .A(\marbiter/_0700_ ), .Z(\wstrb[7] ) );
BUF_X1 \marbiter/_1301_ ( .A(\lsu_wdata[0] ), .Z(\marbiter/_0607_ ) );
BUF_X1 \marbiter/_1302_ ( .A(_351_ ), .Z(\marbiter/_0575_ ) );
BUF_X1 \marbiter/_1303_ ( .A(\marbiter/_0639_ ), .Z(\wdata[0] ) );
BUF_X1 \marbiter/_1304_ ( .A(\lsu_wdata[1] ), .Z(\marbiter/_0618_ ) );
BUF_X1 \marbiter/_1305_ ( .A(_351_ ), .Z(\marbiter/_0586_ ) );
BUF_X1 \marbiter/_1306_ ( .A(\marbiter/_0650_ ), .Z(\wdata[1] ) );
BUF_X1 \marbiter/_1307_ ( .A(\lsu_wdata[2] ), .Z(\marbiter/_0629_ ) );
BUF_X1 \marbiter/_1308_ ( .A(_351_ ), .Z(\marbiter/_0597_ ) );
BUF_X1 \marbiter/_1309_ ( .A(\marbiter/_0661_ ), .Z(\wdata[2] ) );
BUF_X1 \marbiter/_1310_ ( .A(\lsu_wdata[3] ), .Z(\marbiter/_0632_ ) );
BUF_X1 \marbiter/_1311_ ( .A(_351_ ), .Z(\marbiter/_0600_ ) );
BUF_X1 \marbiter/_1312_ ( .A(\marbiter/_0664_ ), .Z(\wdata[3] ) );
BUF_X1 \marbiter/_1313_ ( .A(\lsu_wdata[4] ), .Z(\marbiter/_0633_ ) );
BUF_X1 \marbiter/_1314_ ( .A(_351_ ), .Z(\marbiter/_0601_ ) );
BUF_X1 \marbiter/_1315_ ( .A(\marbiter/_0665_ ), .Z(\wdata[4] ) );
BUF_X1 \marbiter/_1316_ ( .A(\lsu_wdata[5] ), .Z(\marbiter/_0634_ ) );
BUF_X1 \marbiter/_1317_ ( .A(_351_ ), .Z(\marbiter/_0602_ ) );
BUF_X1 \marbiter/_1318_ ( .A(\marbiter/_0666_ ), .Z(\wdata[5] ) );
BUF_X1 \marbiter/_1319_ ( .A(\lsu_wdata[6] ), .Z(\marbiter/_0635_ ) );
BUF_X1 \marbiter/_1320_ ( .A(_351_ ), .Z(\marbiter/_0603_ ) );
BUF_X1 \marbiter/_1321_ ( .A(\marbiter/_0667_ ), .Z(\wdata[6] ) );
BUF_X1 \marbiter/_1322_ ( .A(\lsu_wdata[7] ), .Z(\marbiter/_0636_ ) );
BUF_X1 \marbiter/_1323_ ( .A(_351_ ), .Z(\marbiter/_0604_ ) );
BUF_X1 \marbiter/_1324_ ( .A(\marbiter/_0668_ ), .Z(\wdata[7] ) );
BUF_X1 \marbiter/_1325_ ( .A(\lsu_wdata[8] ), .Z(\marbiter/_0637_ ) );
BUF_X1 \marbiter/_1326_ ( .A(_351_ ), .Z(\marbiter/_0605_ ) );
BUF_X1 \marbiter/_1327_ ( .A(\marbiter/_0669_ ), .Z(\wdata[8] ) );
BUF_X1 \marbiter/_1328_ ( .A(\lsu_wdata[9] ), .Z(\marbiter/_0638_ ) );
BUF_X1 \marbiter/_1329_ ( .A(_351_ ), .Z(\marbiter/_0606_ ) );
BUF_X1 \marbiter/_1330_ ( .A(\marbiter/_0670_ ), .Z(\wdata[9] ) );
BUF_X1 \marbiter/_1331_ ( .A(\lsu_wdata[10] ), .Z(\marbiter/_0608_ ) );
BUF_X1 \marbiter/_1332_ ( .A(_351_ ), .Z(\marbiter/_0576_ ) );
BUF_X1 \marbiter/_1333_ ( .A(\marbiter/_0640_ ), .Z(\wdata[10] ) );
BUF_X1 \marbiter/_1334_ ( .A(\lsu_wdata[11] ), .Z(\marbiter/_0609_ ) );
BUF_X1 \marbiter/_1335_ ( .A(_351_ ), .Z(\marbiter/_0577_ ) );
BUF_X1 \marbiter/_1336_ ( .A(\marbiter/_0641_ ), .Z(\wdata[11] ) );
BUF_X1 \marbiter/_1337_ ( .A(\lsu_wdata[12] ), .Z(\marbiter/_0610_ ) );
BUF_X1 \marbiter/_1338_ ( .A(_351_ ), .Z(\marbiter/_0578_ ) );
BUF_X1 \marbiter/_1339_ ( .A(\marbiter/_0642_ ), .Z(\wdata[12] ) );
BUF_X1 \marbiter/_1340_ ( .A(\lsu_wdata[13] ), .Z(\marbiter/_0611_ ) );
BUF_X1 \marbiter/_1341_ ( .A(_351_ ), .Z(\marbiter/_0579_ ) );
BUF_X1 \marbiter/_1342_ ( .A(\marbiter/_0643_ ), .Z(\wdata[13] ) );
BUF_X1 \marbiter/_1343_ ( .A(\lsu_wdata[14] ), .Z(\marbiter/_0612_ ) );
BUF_X1 \marbiter/_1344_ ( .A(_351_ ), .Z(\marbiter/_0580_ ) );
BUF_X1 \marbiter/_1345_ ( .A(\marbiter/_0644_ ), .Z(\wdata[14] ) );
BUF_X1 \marbiter/_1346_ ( .A(\lsu_wdata[15] ), .Z(\marbiter/_0613_ ) );
BUF_X1 \marbiter/_1347_ ( .A(_351_ ), .Z(\marbiter/_0581_ ) );
BUF_X1 \marbiter/_1348_ ( .A(\marbiter/_0645_ ), .Z(\wdata[15] ) );
BUF_X1 \marbiter/_1349_ ( .A(\lsu_wdata[16] ), .Z(\marbiter/_0614_ ) );
BUF_X1 \marbiter/_1350_ ( .A(_351_ ), .Z(\marbiter/_0582_ ) );
BUF_X1 \marbiter/_1351_ ( .A(\marbiter/_0646_ ), .Z(\wdata[16] ) );
BUF_X1 \marbiter/_1352_ ( .A(\lsu_wdata[17] ), .Z(\marbiter/_0615_ ) );
BUF_X1 \marbiter/_1353_ ( .A(_351_ ), .Z(\marbiter/_0583_ ) );
BUF_X1 \marbiter/_1354_ ( .A(\marbiter/_0647_ ), .Z(\wdata[17] ) );
BUF_X1 \marbiter/_1355_ ( .A(\lsu_wdata[18] ), .Z(\marbiter/_0616_ ) );
BUF_X1 \marbiter/_1356_ ( .A(_351_ ), .Z(\marbiter/_0584_ ) );
BUF_X1 \marbiter/_1357_ ( .A(\marbiter/_0648_ ), .Z(\wdata[18] ) );
BUF_X1 \marbiter/_1358_ ( .A(\lsu_wdata[19] ), .Z(\marbiter/_0617_ ) );
BUF_X1 \marbiter/_1359_ ( .A(_351_ ), .Z(\marbiter/_0585_ ) );
BUF_X1 \marbiter/_1360_ ( .A(\marbiter/_0649_ ), .Z(\wdata[19] ) );
BUF_X1 \marbiter/_1361_ ( .A(\lsu_wdata[20] ), .Z(\marbiter/_0619_ ) );
BUF_X1 \marbiter/_1362_ ( .A(_351_ ), .Z(\marbiter/_0587_ ) );
BUF_X1 \marbiter/_1363_ ( .A(\marbiter/_0651_ ), .Z(\wdata[20] ) );
BUF_X1 \marbiter/_1364_ ( .A(\lsu_wdata[21] ), .Z(\marbiter/_0620_ ) );
BUF_X1 \marbiter/_1365_ ( .A(_351_ ), .Z(\marbiter/_0588_ ) );
BUF_X1 \marbiter/_1366_ ( .A(\marbiter/_0652_ ), .Z(\wdata[21] ) );
BUF_X1 \marbiter/_1367_ ( .A(\lsu_wdata[22] ), .Z(\marbiter/_0621_ ) );
BUF_X1 \marbiter/_1368_ ( .A(_351_ ), .Z(\marbiter/_0589_ ) );
BUF_X1 \marbiter/_1369_ ( .A(\marbiter/_0653_ ), .Z(\wdata[22] ) );
BUF_X1 \marbiter/_1370_ ( .A(\lsu_wdata[23] ), .Z(\marbiter/_0622_ ) );
BUF_X1 \marbiter/_1371_ ( .A(_351_ ), .Z(\marbiter/_0590_ ) );
BUF_X1 \marbiter/_1372_ ( .A(\marbiter/_0654_ ), .Z(\wdata[23] ) );
BUF_X1 \marbiter/_1373_ ( .A(\lsu_wdata[24] ), .Z(\marbiter/_0623_ ) );
BUF_X1 \marbiter/_1374_ ( .A(_351_ ), .Z(\marbiter/_0591_ ) );
BUF_X1 \marbiter/_1375_ ( .A(\marbiter/_0655_ ), .Z(\wdata[24] ) );
BUF_X1 \marbiter/_1376_ ( .A(\lsu_wdata[25] ), .Z(\marbiter/_0624_ ) );
BUF_X1 \marbiter/_1377_ ( .A(_351_ ), .Z(\marbiter/_0592_ ) );
BUF_X1 \marbiter/_1378_ ( .A(\marbiter/_0656_ ), .Z(\wdata[25] ) );
BUF_X1 \marbiter/_1379_ ( .A(\lsu_wdata[26] ), .Z(\marbiter/_0625_ ) );
BUF_X1 \marbiter/_1380_ ( .A(_351_ ), .Z(\marbiter/_0593_ ) );
BUF_X1 \marbiter/_1381_ ( .A(\marbiter/_0657_ ), .Z(\wdata[26] ) );
BUF_X1 \marbiter/_1382_ ( .A(\lsu_wdata[27] ), .Z(\marbiter/_0626_ ) );
BUF_X1 \marbiter/_1383_ ( .A(_351_ ), .Z(\marbiter/_0594_ ) );
BUF_X1 \marbiter/_1384_ ( .A(\marbiter/_0658_ ), .Z(\wdata[27] ) );
BUF_X1 \marbiter/_1385_ ( .A(\lsu_wdata[28] ), .Z(\marbiter/_0627_ ) );
BUF_X1 \marbiter/_1386_ ( .A(_351_ ), .Z(\marbiter/_0595_ ) );
BUF_X1 \marbiter/_1387_ ( .A(\marbiter/_0659_ ), .Z(\wdata[28] ) );
BUF_X1 \marbiter/_1388_ ( .A(\lsu_wdata[29] ), .Z(\marbiter/_0628_ ) );
BUF_X1 \marbiter/_1389_ ( .A(_351_ ), .Z(\marbiter/_0596_ ) );
BUF_X1 \marbiter/_1390_ ( .A(\marbiter/_0660_ ), .Z(\wdata[29] ) );
BUF_X1 \marbiter/_1391_ ( .A(\lsu_wdata[30] ), .Z(\marbiter/_0630_ ) );
BUF_X1 \marbiter/_1392_ ( .A(_351_ ), .Z(\marbiter/_0598_ ) );
BUF_X1 \marbiter/_1393_ ( .A(\marbiter/_0662_ ), .Z(\wdata[30] ) );
BUF_X1 \marbiter/_1394_ ( .A(\lsu_wdata[31] ), .Z(\marbiter/_0631_ ) );
BUF_X1 \marbiter/_1395_ ( .A(_351_ ), .Z(\marbiter/_0599_ ) );
BUF_X1 \marbiter/_1396_ ( .A(\marbiter/_0663_ ), .Z(\wdata[31] ) );
BUF_X1 \marbiter/_1397_ ( .A(\lsu_awaddr[0] ), .Z(\marbiter/_0146_ ) );
BUF_X1 \marbiter/_1398_ ( .A(_351_ ), .Z(\marbiter/_0114_ ) );
BUF_X1 \marbiter/_1399_ ( .A(\marbiter/_0178_ ), .Z(\awaddr[0] ) );
BUF_X1 \marbiter/_1400_ ( .A(\lsu_awaddr[1] ), .Z(\marbiter/_0157_ ) );
BUF_X1 \marbiter/_1401_ ( .A(_351_ ), .Z(\marbiter/_0125_ ) );
BUF_X1 \marbiter/_1402_ ( .A(\marbiter/_0189_ ), .Z(\awaddr[1] ) );
BUF_X1 \marbiter/_1403_ ( .A(\lsu_awaddr[2] ), .Z(\marbiter/_0168_ ) );
BUF_X1 \marbiter/_1404_ ( .A(_351_ ), .Z(\marbiter/_0136_ ) );
BUF_X1 \marbiter/_1405_ ( .A(\marbiter/_0200_ ), .Z(\awaddr[2] ) );
BUF_X1 \marbiter/_1406_ ( .A(\lsu_awaddr[3] ), .Z(\marbiter/_0171_ ) );
BUF_X1 \marbiter/_1407_ ( .A(_351_ ), .Z(\marbiter/_0139_ ) );
BUF_X1 \marbiter/_1408_ ( .A(\marbiter/_0203_ ), .Z(\awaddr[3] ) );
BUF_X1 \marbiter/_1409_ ( .A(\lsu_awaddr[4] ), .Z(\marbiter/_0172_ ) );
BUF_X1 \marbiter/_1410_ ( .A(_351_ ), .Z(\marbiter/_0140_ ) );
BUF_X1 \marbiter/_1411_ ( .A(\marbiter/_0204_ ), .Z(\awaddr[4] ) );
BUF_X1 \marbiter/_1412_ ( .A(\lsu_awaddr[5] ), .Z(\marbiter/_0173_ ) );
BUF_X1 \marbiter/_1413_ ( .A(_351_ ), .Z(\marbiter/_0141_ ) );
BUF_X1 \marbiter/_1414_ ( .A(\marbiter/_0205_ ), .Z(\awaddr[5] ) );
BUF_X1 \marbiter/_1415_ ( .A(\lsu_awaddr[6] ), .Z(\marbiter/_0174_ ) );
BUF_X1 \marbiter/_1416_ ( .A(_351_ ), .Z(\marbiter/_0142_ ) );
BUF_X1 \marbiter/_1417_ ( .A(\marbiter/_0206_ ), .Z(\awaddr[6] ) );
BUF_X1 \marbiter/_1418_ ( .A(\lsu_awaddr[7] ), .Z(\marbiter/_0175_ ) );
BUF_X1 \marbiter/_1419_ ( .A(_351_ ), .Z(\marbiter/_0143_ ) );
BUF_X1 \marbiter/_1420_ ( .A(\marbiter/_0207_ ), .Z(\awaddr[7] ) );
BUF_X1 \marbiter/_1421_ ( .A(\lsu_awaddr[8] ), .Z(\marbiter/_0176_ ) );
BUF_X1 \marbiter/_1422_ ( .A(_351_ ), .Z(\marbiter/_0144_ ) );
BUF_X1 \marbiter/_1423_ ( .A(\marbiter/_0208_ ), .Z(\awaddr[8] ) );
BUF_X1 \marbiter/_1424_ ( .A(\lsu_awaddr[9] ), .Z(\marbiter/_0177_ ) );
BUF_X1 \marbiter/_1425_ ( .A(_351_ ), .Z(\marbiter/_0145_ ) );
BUF_X1 \marbiter/_1426_ ( .A(\marbiter/_0209_ ), .Z(\awaddr[9] ) );
BUF_X1 \marbiter/_1427_ ( .A(\lsu_awaddr[10] ), .Z(\marbiter/_0147_ ) );
BUF_X1 \marbiter/_1428_ ( .A(_351_ ), .Z(\marbiter/_0115_ ) );
BUF_X1 \marbiter/_1429_ ( .A(\marbiter/_0179_ ), .Z(\awaddr[10] ) );
BUF_X1 \marbiter/_1430_ ( .A(\lsu_awaddr[11] ), .Z(\marbiter/_0148_ ) );
BUF_X1 \marbiter/_1431_ ( .A(_351_ ), .Z(\marbiter/_0116_ ) );
BUF_X1 \marbiter/_1432_ ( .A(\marbiter/_0180_ ), .Z(\awaddr[11] ) );
BUF_X1 \marbiter/_1433_ ( .A(\lsu_awaddr[12] ), .Z(\marbiter/_0149_ ) );
BUF_X1 \marbiter/_1434_ ( .A(_351_ ), .Z(\marbiter/_0117_ ) );
BUF_X1 \marbiter/_1435_ ( .A(\marbiter/_0181_ ), .Z(\awaddr[12] ) );
BUF_X1 \marbiter/_1436_ ( .A(\lsu_awaddr[13] ), .Z(\marbiter/_0150_ ) );
BUF_X1 \marbiter/_1437_ ( .A(_351_ ), .Z(\marbiter/_0118_ ) );
BUF_X1 \marbiter/_1438_ ( .A(\marbiter/_0182_ ), .Z(\awaddr[13] ) );
BUF_X1 \marbiter/_1439_ ( .A(\lsu_awaddr[14] ), .Z(\marbiter/_0151_ ) );
BUF_X1 \marbiter/_1440_ ( .A(_351_ ), .Z(\marbiter/_0119_ ) );
BUF_X1 \marbiter/_1441_ ( .A(\marbiter/_0183_ ), .Z(\awaddr[14] ) );
BUF_X1 \marbiter/_1442_ ( .A(\lsu_awaddr[15] ), .Z(\marbiter/_0152_ ) );
BUF_X1 \marbiter/_1443_ ( .A(_351_ ), .Z(\marbiter/_0120_ ) );
BUF_X1 \marbiter/_1444_ ( .A(\marbiter/_0184_ ), .Z(\awaddr[15] ) );
BUF_X1 \marbiter/_1445_ ( .A(\lsu_awaddr[16] ), .Z(\marbiter/_0153_ ) );
BUF_X1 \marbiter/_1446_ ( .A(_351_ ), .Z(\marbiter/_0121_ ) );
BUF_X1 \marbiter/_1447_ ( .A(\marbiter/_0185_ ), .Z(\awaddr[16] ) );
BUF_X1 \marbiter/_1448_ ( .A(\lsu_awaddr[17] ), .Z(\marbiter/_0154_ ) );
BUF_X1 \marbiter/_1449_ ( .A(_351_ ), .Z(\marbiter/_0122_ ) );
BUF_X1 \marbiter/_1450_ ( .A(\marbiter/_0186_ ), .Z(\awaddr[17] ) );
BUF_X1 \marbiter/_1451_ ( .A(\lsu_awaddr[18] ), .Z(\marbiter/_0155_ ) );
BUF_X1 \marbiter/_1452_ ( .A(_351_ ), .Z(\marbiter/_0123_ ) );
BUF_X1 \marbiter/_1453_ ( .A(\marbiter/_0187_ ), .Z(\awaddr[18] ) );
BUF_X1 \marbiter/_1454_ ( .A(\lsu_awaddr[19] ), .Z(\marbiter/_0156_ ) );
BUF_X1 \marbiter/_1455_ ( .A(_351_ ), .Z(\marbiter/_0124_ ) );
BUF_X1 \marbiter/_1456_ ( .A(\marbiter/_0188_ ), .Z(\awaddr[19] ) );
BUF_X1 \marbiter/_1457_ ( .A(\lsu_awaddr[20] ), .Z(\marbiter/_0158_ ) );
BUF_X1 \marbiter/_1458_ ( .A(_351_ ), .Z(\marbiter/_0126_ ) );
BUF_X1 \marbiter/_1459_ ( .A(\marbiter/_0190_ ), .Z(\awaddr[20] ) );
BUF_X1 \marbiter/_1460_ ( .A(\lsu_awaddr[21] ), .Z(\marbiter/_0159_ ) );
BUF_X1 \marbiter/_1461_ ( .A(_351_ ), .Z(\marbiter/_0127_ ) );
BUF_X1 \marbiter/_1462_ ( .A(\marbiter/_0191_ ), .Z(\awaddr[21] ) );
BUF_X1 \marbiter/_1463_ ( .A(\lsu_awaddr[22] ), .Z(\marbiter/_0160_ ) );
BUF_X1 \marbiter/_1464_ ( .A(_351_ ), .Z(\marbiter/_0128_ ) );
BUF_X1 \marbiter/_1465_ ( .A(\marbiter/_0192_ ), .Z(\awaddr[22] ) );
BUF_X1 \marbiter/_1466_ ( .A(\lsu_awaddr[23] ), .Z(\marbiter/_0161_ ) );
BUF_X1 \marbiter/_1467_ ( .A(_351_ ), .Z(\marbiter/_0129_ ) );
BUF_X1 \marbiter/_1468_ ( .A(\marbiter/_0193_ ), .Z(\awaddr[23] ) );
BUF_X1 \marbiter/_1469_ ( .A(\lsu_awaddr[24] ), .Z(\marbiter/_0162_ ) );
BUF_X1 \marbiter/_1470_ ( .A(_351_ ), .Z(\marbiter/_0130_ ) );
BUF_X1 \marbiter/_1471_ ( .A(\marbiter/_0194_ ), .Z(\awaddr[24] ) );
BUF_X1 \marbiter/_1472_ ( .A(\lsu_awaddr[25] ), .Z(\marbiter/_0163_ ) );
BUF_X1 \marbiter/_1473_ ( .A(_351_ ), .Z(\marbiter/_0131_ ) );
BUF_X1 \marbiter/_1474_ ( .A(\marbiter/_0195_ ), .Z(\awaddr[25] ) );
BUF_X1 \marbiter/_1475_ ( .A(\lsu_awaddr[26] ), .Z(\marbiter/_0164_ ) );
BUF_X1 \marbiter/_1476_ ( .A(_351_ ), .Z(\marbiter/_0132_ ) );
BUF_X1 \marbiter/_1477_ ( .A(\marbiter/_0196_ ), .Z(\awaddr[26] ) );
BUF_X1 \marbiter/_1478_ ( .A(\lsu_awaddr[27] ), .Z(\marbiter/_0165_ ) );
BUF_X1 \marbiter/_1479_ ( .A(_351_ ), .Z(\marbiter/_0133_ ) );
BUF_X1 \marbiter/_1480_ ( .A(\marbiter/_0197_ ), .Z(\awaddr[27] ) );
BUF_X1 \marbiter/_1481_ ( .A(\lsu_awaddr[28] ), .Z(\marbiter/_0166_ ) );
BUF_X1 \marbiter/_1482_ ( .A(_351_ ), .Z(\marbiter/_0134_ ) );
BUF_X1 \marbiter/_1483_ ( .A(\marbiter/_0198_ ), .Z(\awaddr[28] ) );
BUF_X1 \marbiter/_1484_ ( .A(\lsu_awaddr[29] ), .Z(\marbiter/_0167_ ) );
BUF_X1 \marbiter/_1485_ ( .A(_351_ ), .Z(\marbiter/_0135_ ) );
BUF_X1 \marbiter/_1486_ ( .A(\marbiter/_0199_ ), .Z(\awaddr[29] ) );
BUF_X1 \marbiter/_1487_ ( .A(\lsu_awaddr[30] ), .Z(\marbiter/_0169_ ) );
BUF_X1 \marbiter/_1488_ ( .A(_351_ ), .Z(\marbiter/_0137_ ) );
BUF_X1 \marbiter/_1489_ ( .A(\marbiter/_0201_ ), .Z(\awaddr[30] ) );
BUF_X1 \marbiter/_1490_ ( .A(\lsu_awaddr[31] ), .Z(\marbiter/_0170_ ) );
BUF_X1 \marbiter/_1491_ ( .A(_351_ ), .Z(\marbiter/_0138_ ) );
BUF_X1 \marbiter/_1492_ ( .A(\marbiter/_0202_ ), .Z(\awaddr[31] ) );
BUF_X1 \marbiter/_1493_ ( .A(lsu_bready ), .Z(\marbiter/_0218_ ) );
BUF_X1 \marbiter/_1494_ ( .A(_351_ ), .Z(\marbiter/_0217_ ) );
BUF_X1 \marbiter/_1495_ ( .A(\marbiter/_0216_ ), .Z(bready ) );
BUF_X1 \marbiter/_1496_ ( .A(\marbiter/_0701_ ), .Z(wvalid ) );
BUF_X1 \marbiter/_1497_ ( .A(\marbiter/_0213_ ), .Z(awvalid ) );
BUF_X1 \marbiter/_1498_ ( .A(\lsu_araddr[0] ), .Z(\marbiter/_0044_ ) );
BUF_X1 \marbiter/_1499_ ( .A(\ifu_araddr[0] ), .Z(\marbiter/_0012_ ) );
BUF_X1 \marbiter/_1500_ ( .A(\marbiter/_0076_ ), .Z(\araddr[0] ) );
BUF_X1 \marbiter/_1501_ ( .A(\lsu_araddr[1] ), .Z(\marbiter/_0055_ ) );
BUF_X1 \marbiter/_1502_ ( .A(\ifu_araddr[1] ), .Z(\marbiter/_0023_ ) );
BUF_X1 \marbiter/_1503_ ( .A(\marbiter/_0087_ ), .Z(\araddr[1] ) );
BUF_X1 \marbiter/_1504_ ( .A(\lsu_araddr[2] ), .Z(\marbiter/_0066_ ) );
BUF_X1 \marbiter/_1505_ ( .A(\ifu_araddr[2] ), .Z(\marbiter/_0034_ ) );
BUF_X1 \marbiter/_1506_ ( .A(\marbiter/_0098_ ), .Z(\araddr[2] ) );
BUF_X1 \marbiter/_1507_ ( .A(\lsu_araddr[3] ), .Z(\marbiter/_0069_ ) );
BUF_X1 \marbiter/_1508_ ( .A(\ifu_araddr[3] ), .Z(\marbiter/_0037_ ) );
BUF_X1 \marbiter/_1509_ ( .A(\marbiter/_0101_ ), .Z(\araddr[3] ) );
BUF_X1 \marbiter/_1510_ ( .A(\lsu_araddr[4] ), .Z(\marbiter/_0070_ ) );
BUF_X1 \marbiter/_1511_ ( .A(\ifu_araddr[4] ), .Z(\marbiter/_0038_ ) );
BUF_X1 \marbiter/_1512_ ( .A(\marbiter/_0102_ ), .Z(\araddr[4] ) );
BUF_X1 \marbiter/_1513_ ( .A(\lsu_araddr[5] ), .Z(\marbiter/_0071_ ) );
BUF_X1 \marbiter/_1514_ ( .A(\ifu_araddr[5] ), .Z(\marbiter/_0039_ ) );
BUF_X1 \marbiter/_1515_ ( .A(\marbiter/_0103_ ), .Z(\araddr[5] ) );
BUF_X1 \marbiter/_1516_ ( .A(\lsu_araddr[6] ), .Z(\marbiter/_0072_ ) );
BUF_X1 \marbiter/_1517_ ( .A(\ifu_araddr[6] ), .Z(\marbiter/_0040_ ) );
BUF_X1 \marbiter/_1518_ ( .A(\marbiter/_0104_ ), .Z(\araddr[6] ) );
BUF_X1 \marbiter/_1519_ ( .A(\lsu_araddr[7] ), .Z(\marbiter/_0073_ ) );
BUF_X1 \marbiter/_1520_ ( .A(\ifu_araddr[7] ), .Z(\marbiter/_0041_ ) );
BUF_X1 \marbiter/_1521_ ( .A(\marbiter/_0105_ ), .Z(\araddr[7] ) );
BUF_X1 \marbiter/_1522_ ( .A(\lsu_araddr[8] ), .Z(\marbiter/_0074_ ) );
BUF_X1 \marbiter/_1523_ ( .A(\ifu_araddr[8] ), .Z(\marbiter/_0042_ ) );
BUF_X1 \marbiter/_1524_ ( .A(\marbiter/_0106_ ), .Z(\araddr[8] ) );
BUF_X1 \marbiter/_1525_ ( .A(\lsu_araddr[9] ), .Z(\marbiter/_0075_ ) );
BUF_X1 \marbiter/_1526_ ( .A(\ifu_araddr[9] ), .Z(\marbiter/_0043_ ) );
BUF_X1 \marbiter/_1527_ ( .A(\marbiter/_0107_ ), .Z(\araddr[9] ) );
BUF_X1 \marbiter/_1528_ ( .A(\lsu_araddr[10] ), .Z(\marbiter/_0045_ ) );
BUF_X1 \marbiter/_1529_ ( .A(\ifu_araddr[10] ), .Z(\marbiter/_0013_ ) );
BUF_X1 \marbiter/_1530_ ( .A(\marbiter/_0077_ ), .Z(\araddr[10] ) );
BUF_X1 \marbiter/_1531_ ( .A(\lsu_araddr[11] ), .Z(\marbiter/_0046_ ) );
BUF_X1 \marbiter/_1532_ ( .A(\ifu_araddr[11] ), .Z(\marbiter/_0014_ ) );
BUF_X1 \marbiter/_1533_ ( .A(\marbiter/_0078_ ), .Z(\araddr[11] ) );
BUF_X1 \marbiter/_1534_ ( .A(\lsu_araddr[12] ), .Z(\marbiter/_0047_ ) );
BUF_X1 \marbiter/_1535_ ( .A(\ifu_araddr[12] ), .Z(\marbiter/_0015_ ) );
BUF_X1 \marbiter/_1536_ ( .A(\marbiter/_0079_ ), .Z(\araddr[12] ) );
BUF_X1 \marbiter/_1537_ ( .A(\lsu_araddr[13] ), .Z(\marbiter/_0048_ ) );
BUF_X1 \marbiter/_1538_ ( .A(\ifu_araddr[13] ), .Z(\marbiter/_0016_ ) );
BUF_X1 \marbiter/_1539_ ( .A(\marbiter/_0080_ ), .Z(\araddr[13] ) );
BUF_X1 \marbiter/_1540_ ( .A(\lsu_araddr[14] ), .Z(\marbiter/_0049_ ) );
BUF_X1 \marbiter/_1541_ ( .A(\ifu_araddr[14] ), .Z(\marbiter/_0017_ ) );
BUF_X1 \marbiter/_1542_ ( .A(\marbiter/_0081_ ), .Z(\araddr[14] ) );
BUF_X1 \marbiter/_1543_ ( .A(\lsu_araddr[15] ), .Z(\marbiter/_0050_ ) );
BUF_X1 \marbiter/_1544_ ( .A(\ifu_araddr[15] ), .Z(\marbiter/_0018_ ) );
BUF_X1 \marbiter/_1545_ ( .A(\marbiter/_0082_ ), .Z(\araddr[15] ) );
BUF_X1 \marbiter/_1546_ ( .A(\lsu_araddr[16] ), .Z(\marbiter/_0051_ ) );
BUF_X1 \marbiter/_1547_ ( .A(\ifu_araddr[16] ), .Z(\marbiter/_0019_ ) );
BUF_X1 \marbiter/_1548_ ( .A(\marbiter/_0083_ ), .Z(\araddr[16] ) );
BUF_X1 \marbiter/_1549_ ( .A(\lsu_araddr[17] ), .Z(\marbiter/_0052_ ) );
BUF_X1 \marbiter/_1550_ ( .A(\ifu_araddr[17] ), .Z(\marbiter/_0020_ ) );
BUF_X1 \marbiter/_1551_ ( .A(\marbiter/_0084_ ), .Z(\araddr[17] ) );
BUF_X1 \marbiter/_1552_ ( .A(\lsu_araddr[18] ), .Z(\marbiter/_0053_ ) );
BUF_X1 \marbiter/_1553_ ( .A(\ifu_araddr[18] ), .Z(\marbiter/_0021_ ) );
BUF_X1 \marbiter/_1554_ ( .A(\marbiter/_0085_ ), .Z(\araddr[18] ) );
BUF_X1 \marbiter/_1555_ ( .A(\lsu_araddr[19] ), .Z(\marbiter/_0054_ ) );
BUF_X1 \marbiter/_1556_ ( .A(\ifu_araddr[19] ), .Z(\marbiter/_0022_ ) );
BUF_X1 \marbiter/_1557_ ( .A(\marbiter/_0086_ ), .Z(\araddr[19] ) );
BUF_X1 \marbiter/_1558_ ( .A(\lsu_araddr[20] ), .Z(\marbiter/_0056_ ) );
BUF_X1 \marbiter/_1559_ ( .A(\ifu_araddr[20] ), .Z(\marbiter/_0024_ ) );
BUF_X1 \marbiter/_1560_ ( .A(\marbiter/_0088_ ), .Z(\araddr[20] ) );
BUF_X1 \marbiter/_1561_ ( .A(\lsu_araddr[21] ), .Z(\marbiter/_0057_ ) );
BUF_X1 \marbiter/_1562_ ( .A(\ifu_araddr[21] ), .Z(\marbiter/_0025_ ) );
BUF_X1 \marbiter/_1563_ ( .A(\marbiter/_0089_ ), .Z(\araddr[21] ) );
BUF_X1 \marbiter/_1564_ ( .A(\lsu_araddr[22] ), .Z(\marbiter/_0058_ ) );
BUF_X1 \marbiter/_1565_ ( .A(\ifu_araddr[22] ), .Z(\marbiter/_0026_ ) );
BUF_X1 \marbiter/_1566_ ( .A(\marbiter/_0090_ ), .Z(\araddr[22] ) );
BUF_X1 \marbiter/_1567_ ( .A(\lsu_araddr[23] ), .Z(\marbiter/_0059_ ) );
BUF_X1 \marbiter/_1568_ ( .A(\ifu_araddr[23] ), .Z(\marbiter/_0027_ ) );
BUF_X1 \marbiter/_1569_ ( .A(\marbiter/_0091_ ), .Z(\araddr[23] ) );
BUF_X1 \marbiter/_1570_ ( .A(\lsu_araddr[24] ), .Z(\marbiter/_0060_ ) );
BUF_X1 \marbiter/_1571_ ( .A(\ifu_araddr[24] ), .Z(\marbiter/_0028_ ) );
BUF_X1 \marbiter/_1572_ ( .A(\marbiter/_0092_ ), .Z(\araddr[24] ) );
BUF_X1 \marbiter/_1573_ ( .A(\lsu_araddr[25] ), .Z(\marbiter/_0061_ ) );
BUF_X1 \marbiter/_1574_ ( .A(\ifu_araddr[25] ), .Z(\marbiter/_0029_ ) );
BUF_X1 \marbiter/_1575_ ( .A(\marbiter/_0093_ ), .Z(\araddr[25] ) );
BUF_X1 \marbiter/_1576_ ( .A(\lsu_araddr[26] ), .Z(\marbiter/_0062_ ) );
BUF_X1 \marbiter/_1577_ ( .A(\ifu_araddr[26] ), .Z(\marbiter/_0030_ ) );
BUF_X1 \marbiter/_1578_ ( .A(\marbiter/_0094_ ), .Z(\araddr[26] ) );
BUF_X1 \marbiter/_1579_ ( .A(\lsu_araddr[27] ), .Z(\marbiter/_0063_ ) );
BUF_X1 \marbiter/_1580_ ( .A(\ifu_araddr[27] ), .Z(\marbiter/_0031_ ) );
BUF_X1 \marbiter/_1581_ ( .A(\marbiter/_0095_ ), .Z(\araddr[27] ) );
BUF_X1 \marbiter/_1582_ ( .A(\lsu_araddr[28] ), .Z(\marbiter/_0064_ ) );
BUF_X1 \marbiter/_1583_ ( .A(\ifu_araddr[28] ), .Z(\marbiter/_0032_ ) );
BUF_X1 \marbiter/_1584_ ( .A(\marbiter/_0096_ ), .Z(\araddr[28] ) );
BUF_X1 \marbiter/_1585_ ( .A(\lsu_araddr[29] ), .Z(\marbiter/_0065_ ) );
BUF_X1 \marbiter/_1586_ ( .A(\ifu_araddr[29] ), .Z(\marbiter/_0033_ ) );
BUF_X1 \marbiter/_1587_ ( .A(\marbiter/_0097_ ), .Z(\araddr[29] ) );
BUF_X1 \marbiter/_1588_ ( .A(\lsu_araddr[30] ), .Z(\marbiter/_0067_ ) );
BUF_X1 \marbiter/_1589_ ( .A(\ifu_araddr[30] ), .Z(\marbiter/_0035_ ) );
BUF_X1 \marbiter/_1590_ ( .A(\marbiter/_0099_ ), .Z(\araddr[30] ) );
BUF_X1 \marbiter/_1591_ ( .A(\lsu_araddr[31] ), .Z(\marbiter/_0068_ ) );
BUF_X1 \marbiter/_1592_ ( .A(\ifu_araddr[31] ), .Z(\marbiter/_0036_ ) );
BUF_X1 \marbiter/_1593_ ( .A(\marbiter/_0100_ ), .Z(\araddr[31] ) );
BUF_X1 \marbiter/_1594_ ( .A(lsu_rready ), .Z(\marbiter/_0564_ ) );
BUF_X1 \marbiter/_1595_ ( .A(ifu_rready ), .Z(\marbiter/_0563_ ) );
BUF_X1 \marbiter/_1596_ ( .A(\marbiter/_0562_ ), .Z(rready ) );
BUF_X1 \marbiter/_1597_ ( .A(\marbiter/_0111_ ), .Z(arvalid ) );
BUF_X1 \marbiter/_1598_ ( .A(arready ), .Z(\marbiter/_0108_ ) );
BUF_X1 \marbiter/_1599_ ( .A(\marbiter/_0109_ ), .Z(ifu_arready ) );
BUF_X1 \marbiter/_1600_ ( .A(\marbiter/_0573_ ), .Z(ifu_rvalid ) );
BUF_X1 \marbiter/_1601_ ( .A(\marbiter/_0110_ ), .Z(lsu_arready ) );
BUF_X1 \marbiter/_1602_ ( .A(\marbiter/_0574_ ), .Z(lsu_rvalid ) );
BUF_X1 \marbiter/_1603_ ( .A(awready ), .Z(\marbiter/_0210_ ) );
BUF_X1 \marbiter/_1604_ ( .A(\marbiter/_0211_ ), .Z(ifu_awready ) );
BUF_X1 \marbiter/_1605_ ( .A(\marbiter/_0672_ ), .Z(ifu_wready ) );
BUF_X1 \marbiter/_1606_ ( .A(bvalid ), .Z(\marbiter/_0225_ ) );
BUF_X1 \marbiter/_1607_ ( .A(\marbiter/_0226_ ), .Z(ifu_bvalid ) );
BUF_X1 \marbiter/_1608_ ( .A(\marbiter/_0212_ ), .Z(lsu_awready ) );
BUF_X1 \marbiter/_1609_ ( .A(\marbiter/_0673_ ), .Z(lsu_wready ) );
BUF_X1 \marbiter/_1610_ ( .A(\marbiter/_0227_ ), .Z(lsu_bvalid ) );
AND2_X1 \mcsr/_1155_ ( .A1(\mcsr/_0267_ ), .A2(\mcsr/_0266_ ), .ZN(\mcsr/_0334_ ) );
NOR2_X1 \mcsr/_1156_ ( .A1(\mcsr/_0258_ ), .A2(\mcsr/_0257_ ), .ZN(\mcsr/_0335_ ) );
AND2_X2 \mcsr/_1157_ ( .A1(\mcsr/_0334_ ), .A2(\mcsr/_0335_ ), .ZN(\mcsr/_0336_ ) );
INV_X1 \mcsr/_1158_ ( .A(\mcsr/_0264_ ), .ZN(\mcsr/_0337_ ) );
NOR4_X4 \mcsr/_1159_ ( .A1(\mcsr/_0337_ ), .A2(\mcsr/_0261_ ), .A3(\mcsr/_0260_ ), .A4(\mcsr/_0265_ ), .ZN(\mcsr/_0338_ ) );
AND2_X4 \mcsr/_1160_ ( .A1(\mcsr/_0336_ ), .A2(\mcsr/_0338_ ), .ZN(\mcsr/_0339_ ) );
INV_X2 \mcsr/_1161_ ( .A(\mcsr/_0259_ ), .ZN(\mcsr/_0340_ ) );
NOR4_X4 \mcsr/_1162_ ( .A1(\mcsr/_0340_ ), .A2(\mcsr/_0256_ ), .A3(\mcsr/_0263_ ), .A4(\mcsr/_0262_ ), .ZN(\mcsr/_0341_ ) );
AND2_X4 \mcsr/_1163_ ( .A1(\mcsr/_0339_ ), .A2(\mcsr/_0341_ ), .ZN(\mcsr/_0342_ ) );
NOR2_X1 \mcsr/_1164_ ( .A1(\mcsr/_0263_ ), .A2(\mcsr/_0262_ ), .ZN(\mcsr/_0343_ ) );
AND3_X1 \mcsr/_1165_ ( .A1(\mcsr/_0343_ ), .A2(\mcsr/_0340_ ), .A3(\mcsr/_0256_ ), .ZN(\mcsr/_0344_ ) );
AND3_X4 \mcsr/_1166_ ( .A1(\mcsr/_0344_ ), .A2(\mcsr/_0336_ ), .A3(\mcsr/_0338_ ), .ZN(\mcsr/_0345_ ) );
NOR2_X4 \mcsr/_1167_ ( .A1(\mcsr/_0342_ ), .A2(\mcsr/_0345_ ), .ZN(\mcsr/_0346_ ) );
NOR2_X1 \mcsr/_1168_ ( .A1(\mcsr/_0261_ ), .A2(\mcsr/_0265_ ), .ZN(\mcsr/_0347_ ) );
AND3_X1 \mcsr/_1169_ ( .A1(\mcsr/_0347_ ), .A2(\mcsr/_0260_ ), .A3(\mcsr/_0337_ ), .ZN(\mcsr/_0348_ ) );
AND2_X1 \mcsr/_1170_ ( .A1(\mcsr/_0348_ ), .A2(\mcsr/_0344_ ), .ZN(\mcsr/_0349_ ) );
AND2_X1 \mcsr/_1171_ ( .A1(\mcsr/_0349_ ), .A2(\mcsr/_0336_ ), .ZN(\mcsr/_0350_ ) );
INV_X1 \mcsr/_1172_ ( .A(\mcsr/_0350_ ), .ZN(\mcsr/_0351_ ) );
AND2_X2 \mcsr/_1173_ ( .A1(\mcsr/_0346_ ), .A2(\mcsr/_0351_ ), .ZN(\mcsr/_0352_ ) );
INV_X1 \mcsr/_1174_ ( .A(\mcsr/_0224_ ), .ZN(\mcsr/_0353_ ) );
INV_X1 \mcsr/_1175_ ( .A(\mcsr/_0343_ ), .ZN(\mcsr/_0354_ ) );
NOR3_X1 \mcsr/_1176_ ( .A1(\mcsr/_0354_ ), .A2(\mcsr/_0265_ ), .A3(\mcsr/_0337_ ), .ZN(\mcsr/_0355_ ) );
NOR4_X1 \mcsr/_1177_ ( .A1(\mcsr/_0340_ ), .A2(\mcsr/_0256_ ), .A3(\mcsr/_0261_ ), .A4(\mcsr/_0260_ ), .ZN(\mcsr/_0356_ ) );
AND3_X1 \mcsr/_1178_ ( .A1(\mcsr/_0355_ ), .A2(\mcsr/_0336_ ), .A3(\mcsr/_0356_ ), .ZN(\mcsr/_0357_ ) );
INV_X1 \mcsr/_1179_ ( .A(\mcsr/_0357_ ), .ZN(\mcsr/_0358_ ) );
AOI21_X1 \mcsr/_1180_ ( .A(\mcsr/_0353_ ), .B1(\mcsr/_0351_ ), .B2(\mcsr/_0358_ ), .ZN(\mcsr/_0359_ ) );
NOR2_X1 \mcsr/_1181_ ( .A1(\mcsr/_0350_ ), .A2(\mcsr/_0357_ ), .ZN(\mcsr/_0360_ ) );
AOI211_X2 \mcsr/_1182_ ( .A(\mcsr/_0346_ ), .B(\mcsr/_0359_ ), .C1(\mcsr/_0192_ ), .C2(\mcsr/_0360_ ), .ZN(\mcsr/_0361_ ) );
NOR2_X1 \mcsr/_1183_ ( .A1(\mcsr/_0350_ ), .A2(\mcsr/_0342_ ), .ZN(\mcsr/_0362_ ) );
OAI22_X1 \mcsr/_1184_ ( .A1(\mcsr/_0362_ ), .A2(\mcsr/_0160_ ), .B1(\mcsr/_0128_ ), .B2(\mcsr/_0350_ ), .ZN(\mcsr/_0363_ ) );
AOI211_X2 \mcsr/_1185_ ( .A(\mcsr/_0352_ ), .B(\mcsr/_0361_ ), .C1(\mcsr/_0346_ ), .C2(\mcsr/_0363_ ), .ZN(\mcsr/_0802_ ) );
BUF_X4 \mcsr/_1186_ ( .A(\mcsr/_0352_ ), .Z(\mcsr/_0364_ ) );
INV_X8 \mcsr/_1187_ ( .A(\mcsr/_0342_ ), .ZN(\mcsr/_0365_ ) );
BUF_X4 \mcsr/_1188_ ( .A(\mcsr/_0365_ ), .Z(\mcsr/_0366_ ) );
INV_X1 \mcsr/_1189_ ( .A(\mcsr/_0345_ ), .ZN(\mcsr/_0367_ ) );
BUF_X4 \mcsr/_1190_ ( .A(\mcsr/_0367_ ), .Z(\mcsr/_0368_ ) );
AND3_X2 \mcsr/_1191_ ( .A1(\mcsr/_0348_ ), .A2(\mcsr/_0344_ ), .A3(\mcsr/_0336_ ), .ZN(\mcsr/_0369_ ) );
INV_X2 \mcsr/_1192_ ( .A(\mcsr/_0369_ ), .ZN(\mcsr/_0370_ ) );
BUF_X4 \mcsr/_1193_ ( .A(\mcsr/_0370_ ), .Z(\mcsr/_0371_ ) );
OAI211_X2 \mcsr/_1194_ ( .A(\mcsr/_0366_ ), .B(\mcsr/_0368_ ), .C1(\mcsr/_0171_ ), .C2(\mcsr/_0371_ ), .ZN(\mcsr/_0372_ ) );
INV_X1 \mcsr/_1195_ ( .A(\mcsr/_0372_ ), .ZN(\mcsr/_0373_ ) );
NOR2_X4 \mcsr/_1196_ ( .A1(\mcsr/_0342_ ), .A2(\mcsr/_0369_ ), .ZN(\mcsr/_0374_ ) );
BUF_X8 \mcsr/_1197_ ( .A(\mcsr/_0374_ ), .Z(\mcsr/_0375_ ) );
INV_X4 \mcsr/_1198_ ( .A(\mcsr/_0375_ ), .ZN(\mcsr/_0376_ ) );
BUF_X4 \mcsr/_1199_ ( .A(\mcsr/_0376_ ), .Z(\mcsr/_0377_ ) );
OAI21_X1 \mcsr/_1200_ ( .A(\mcsr/_0373_ ), .B1(\mcsr/_0139_ ), .B2(\mcsr/_0377_ ), .ZN(\mcsr/_0378_ ) );
INV_X1 \mcsr/_1201_ ( .A(\mcsr/_0346_ ), .ZN(\mcsr/_0379_ ) );
INV_X1 \mcsr/_1202_ ( .A(\mcsr/_0235_ ), .ZN(\mcsr/_0380_ ) );
OAI21_X1 \mcsr/_1203_ ( .A(\mcsr/_0380_ ), .B1(\mcsr/_0342_ ), .B2(\mcsr/_0369_ ), .ZN(\mcsr/_0381_ ) );
OAI211_X2 \mcsr/_1204_ ( .A(\mcsr/_0379_ ), .B(\mcsr/_0381_ ), .C1(\mcsr/_0376_ ), .C2(\mcsr/_0203_ ), .ZN(\mcsr/_0382_ ) );
AOI21_X1 \mcsr/_1205_ ( .A(\mcsr/_0364_ ), .B1(\mcsr/_0378_ ), .B2(\mcsr/_0382_ ), .ZN(\mcsr/_0813_ ) );
OAI211_X2 \mcsr/_1206_ ( .A(\mcsr/_0366_ ), .B(\mcsr/_0368_ ), .C1(\mcsr/_0182_ ), .C2(\mcsr/_0371_ ), .ZN(\mcsr/_0383_ ) );
INV_X1 \mcsr/_1207_ ( .A(\mcsr/_0383_ ), .ZN(\mcsr/_0384_ ) );
OAI21_X1 \mcsr/_1208_ ( .A(\mcsr/_0384_ ), .B1(\mcsr/_0150_ ), .B2(\mcsr/_0377_ ), .ZN(\mcsr/_0385_ ) );
BUF_X8 \mcsr/_1209_ ( .A(\mcsr/_0375_ ), .Z(\mcsr/_0386_ ) );
OR2_X1 \mcsr/_1210_ ( .A1(\mcsr/_0386_ ), .A2(\mcsr/_0246_ ), .ZN(\mcsr/_0387_ ) );
BUF_X4 \mcsr/_1211_ ( .A(\mcsr/_0375_ ), .Z(\mcsr/_0388_ ) );
INV_X1 \mcsr/_1212_ ( .A(\mcsr/_0214_ ), .ZN(\mcsr/_0389_ ) );
BUF_X32 \mcsr/_1213_ ( .A(\mcsr/_0365_ ), .Z(\mcsr/_0390_ ) );
BUF_X32 \mcsr/_1214_ ( .A(\mcsr/_0390_ ), .Z(\mcsr/_0391_ ) );
BUF_X8 \mcsr/_1215_ ( .A(\mcsr/_0367_ ), .Z(\mcsr/_0392_ ) );
BUF_X16 \mcsr/_1216_ ( .A(\mcsr/_0392_ ), .Z(\mcsr/_0393_ ) );
AOI22_X2 \mcsr/_1217_ ( .A1(\mcsr/_0388_ ), .A2(\mcsr/_0389_ ), .B1(\mcsr/_0391_ ), .B2(\mcsr/_0393_ ), .ZN(\mcsr/_0394_ ) );
NAND2_X1 \mcsr/_1218_ ( .A1(\mcsr/_0387_ ), .A2(\mcsr/_0394_ ), .ZN(\mcsr/_0395_ ) );
AOI21_X1 \mcsr/_1219_ ( .A(\mcsr/_0364_ ), .B1(\mcsr/_0385_ ), .B2(\mcsr/_0395_ ), .ZN(\mcsr/_0824_ ) );
OAI211_X2 \mcsr/_1220_ ( .A(\mcsr/_0366_ ), .B(\mcsr/_0368_ ), .C1(\mcsr/_0185_ ), .C2(\mcsr/_0371_ ), .ZN(\mcsr/_0396_ ) );
INV_X1 \mcsr/_1221_ ( .A(\mcsr/_0396_ ), .ZN(\mcsr/_0397_ ) );
OAI21_X1 \mcsr/_1222_ ( .A(\mcsr/_0397_ ), .B1(\mcsr/_0153_ ), .B2(\mcsr/_0377_ ), .ZN(\mcsr/_0398_ ) );
INV_X1 \mcsr/_1223_ ( .A(\mcsr/_0249_ ), .ZN(\mcsr/_0399_ ) );
OAI21_X1 \mcsr/_1224_ ( .A(\mcsr/_0399_ ), .B1(\mcsr/_0342_ ), .B2(\mcsr/_0369_ ), .ZN(\mcsr/_0400_ ) );
OAI211_X2 \mcsr/_1225_ ( .A(\mcsr/_0379_ ), .B(\mcsr/_0400_ ), .C1(\mcsr/_0376_ ), .C2(\mcsr/_0217_ ), .ZN(\mcsr/_0401_ ) );
AOI21_X1 \mcsr/_1226_ ( .A(\mcsr/_0364_ ), .B1(\mcsr/_0398_ ), .B2(\mcsr/_0401_ ), .ZN(\mcsr/_0827_ ) );
BUF_X8 \mcsr/_1227_ ( .A(\mcsr/_0390_ ), .Z(\mcsr/_0402_ ) );
BUF_X8 \mcsr/_1228_ ( .A(\mcsr/_0392_ ), .Z(\mcsr/_0403_ ) );
OAI211_X2 \mcsr/_1229_ ( .A(\mcsr/_0402_ ), .B(\mcsr/_0403_ ), .C1(\mcsr/_0186_ ), .C2(\mcsr/_0371_ ), .ZN(\mcsr/_0404_ ) );
INV_X1 \mcsr/_1230_ ( .A(\mcsr/_0404_ ), .ZN(\mcsr/_0405_ ) );
OAI21_X1 \mcsr/_1231_ ( .A(\mcsr/_0405_ ), .B1(\mcsr/_0154_ ), .B2(\mcsr/_0377_ ), .ZN(\mcsr/_0406_ ) );
OR2_X1 \mcsr/_1232_ ( .A1(\mcsr/_0386_ ), .A2(\mcsr/_0250_ ), .ZN(\mcsr/_0407_ ) );
INV_X1 \mcsr/_1233_ ( .A(\mcsr/_0218_ ), .ZN(\mcsr/_0408_ ) );
AOI22_X2 \mcsr/_1234_ ( .A1(\mcsr/_0388_ ), .A2(\mcsr/_0408_ ), .B1(\mcsr/_0391_ ), .B2(\mcsr/_0393_ ), .ZN(\mcsr/_0409_ ) );
NAND2_X1 \mcsr/_1235_ ( .A1(\mcsr/_0407_ ), .A2(\mcsr/_0409_ ), .ZN(\mcsr/_0410_ ) );
AOI21_X1 \mcsr/_1236_ ( .A(\mcsr/_0364_ ), .B1(\mcsr/_0406_ ), .B2(\mcsr/_0410_ ), .ZN(\mcsr/_0828_ ) );
OAI211_X2 \mcsr/_1237_ ( .A(\mcsr/_0402_ ), .B(\mcsr/_0403_ ), .C1(\mcsr/_0187_ ), .C2(\mcsr/_0371_ ), .ZN(\mcsr/_0411_ ) );
INV_X1 \mcsr/_1238_ ( .A(\mcsr/_0411_ ), .ZN(\mcsr/_0412_ ) );
OAI21_X1 \mcsr/_1239_ ( .A(\mcsr/_0412_ ), .B1(\mcsr/_0155_ ), .B2(\mcsr/_0377_ ), .ZN(\mcsr/_0413_ ) );
OR2_X1 \mcsr/_1240_ ( .A1(\mcsr/_0386_ ), .A2(\mcsr/_0251_ ), .ZN(\mcsr/_0414_ ) );
INV_X1 \mcsr/_1241_ ( .A(\mcsr/_0219_ ), .ZN(\mcsr/_0415_ ) );
AOI22_X2 \mcsr/_1242_ ( .A1(\mcsr/_0388_ ), .A2(\mcsr/_0415_ ), .B1(\mcsr/_0391_ ), .B2(\mcsr/_0393_ ), .ZN(\mcsr/_0416_ ) );
NAND2_X1 \mcsr/_1243_ ( .A1(\mcsr/_0414_ ), .A2(\mcsr/_0416_ ), .ZN(\mcsr/_0417_ ) );
AOI21_X1 \mcsr/_1244_ ( .A(\mcsr/_0364_ ), .B1(\mcsr/_0413_ ), .B2(\mcsr/_0417_ ), .ZN(\mcsr/_0829_ ) );
OAI211_X2 \mcsr/_1245_ ( .A(\mcsr/_0402_ ), .B(\mcsr/_0403_ ), .C1(\mcsr/_0188_ ), .C2(\mcsr/_0371_ ), .ZN(\mcsr/_0418_ ) );
INV_X1 \mcsr/_1246_ ( .A(\mcsr/_0418_ ), .ZN(\mcsr/_0419_ ) );
OAI21_X1 \mcsr/_1247_ ( .A(\mcsr/_0419_ ), .B1(\mcsr/_0156_ ), .B2(\mcsr/_0377_ ), .ZN(\mcsr/_0420_ ) );
CLKBUF_X2 \mcsr/_1248_ ( .A(\mcsr/_0374_ ), .Z(\mcsr/_0421_ ) );
OR2_X1 \mcsr/_1249_ ( .A1(\mcsr/_0421_ ), .A2(\mcsr/_0252_ ), .ZN(\mcsr/_0422_ ) );
INV_X1 \mcsr/_1250_ ( .A(\mcsr/_0220_ ), .ZN(\mcsr/_0423_ ) );
AOI22_X2 \mcsr/_1251_ ( .A1(\mcsr/_0388_ ), .A2(\mcsr/_0423_ ), .B1(\mcsr/_0391_ ), .B2(\mcsr/_0393_ ), .ZN(\mcsr/_0424_ ) );
NAND2_X1 \mcsr/_1252_ ( .A1(\mcsr/_0422_ ), .A2(\mcsr/_0424_ ), .ZN(\mcsr/_0425_ ) );
AOI21_X1 \mcsr/_1253_ ( .A(\mcsr/_0364_ ), .B1(\mcsr/_0420_ ), .B2(\mcsr/_0425_ ), .ZN(\mcsr/_0830_ ) );
OAI211_X2 \mcsr/_1254_ ( .A(\mcsr/_0402_ ), .B(\mcsr/_0403_ ), .C1(\mcsr/_0189_ ), .C2(\mcsr/_0371_ ), .ZN(\mcsr/_0426_ ) );
INV_X1 \mcsr/_1255_ ( .A(\mcsr/_0426_ ), .ZN(\mcsr/_0427_ ) );
OAI21_X1 \mcsr/_1256_ ( .A(\mcsr/_0427_ ), .B1(\mcsr/_0157_ ), .B2(\mcsr/_0377_ ), .ZN(\mcsr/_0428_ ) );
OR2_X1 \mcsr/_1257_ ( .A1(\mcsr/_0421_ ), .A2(\mcsr/_0253_ ), .ZN(\mcsr/_0429_ ) );
INV_X1 \mcsr/_1258_ ( .A(\mcsr/_0221_ ), .ZN(\mcsr/_0430_ ) );
AOI22_X2 \mcsr/_1259_ ( .A1(\mcsr/_0388_ ), .A2(\mcsr/_0430_ ), .B1(\mcsr/_0391_ ), .B2(\mcsr/_0393_ ), .ZN(\mcsr/_0431_ ) );
NAND2_X1 \mcsr/_1260_ ( .A1(\mcsr/_0429_ ), .A2(\mcsr/_0431_ ), .ZN(\mcsr/_0432_ ) );
AOI21_X1 \mcsr/_1261_ ( .A(\mcsr/_0364_ ), .B1(\mcsr/_0428_ ), .B2(\mcsr/_0432_ ), .ZN(\mcsr/_0831_ ) );
OAI211_X2 \mcsr/_1262_ ( .A(\mcsr/_0402_ ), .B(\mcsr/_0403_ ), .C1(\mcsr/_0190_ ), .C2(\mcsr/_0371_ ), .ZN(\mcsr/_0433_ ) );
INV_X1 \mcsr/_1263_ ( .A(\mcsr/_0433_ ), .ZN(\mcsr/_0434_ ) );
OAI21_X1 \mcsr/_1264_ ( .A(\mcsr/_0434_ ), .B1(\mcsr/_0158_ ), .B2(\mcsr/_0377_ ), .ZN(\mcsr/_0435_ ) );
OR2_X1 \mcsr/_1265_ ( .A1(\mcsr/_0421_ ), .A2(\mcsr/_0254_ ), .ZN(\mcsr/_0436_ ) );
INV_X1 \mcsr/_1266_ ( .A(\mcsr/_0222_ ), .ZN(\mcsr/_0437_ ) );
AOI22_X2 \mcsr/_1267_ ( .A1(\mcsr/_0388_ ), .A2(\mcsr/_0437_ ), .B1(\mcsr/_0391_ ), .B2(\mcsr/_0393_ ), .ZN(\mcsr/_0438_ ) );
NAND2_X1 \mcsr/_1268_ ( .A1(\mcsr/_0436_ ), .A2(\mcsr/_0438_ ), .ZN(\mcsr/_0439_ ) );
AOI21_X1 \mcsr/_1269_ ( .A(\mcsr/_0364_ ), .B1(\mcsr/_0435_ ), .B2(\mcsr/_0439_ ), .ZN(\mcsr/_0832_ ) );
BUF_X8 \mcsr/_1270_ ( .A(\mcsr/_0370_ ), .Z(\mcsr/_0440_ ) );
OAI211_X2 \mcsr/_1271_ ( .A(\mcsr/_0402_ ), .B(\mcsr/_0403_ ), .C1(\mcsr/_0191_ ), .C2(\mcsr/_0440_ ), .ZN(\mcsr/_0441_ ) );
INV_X1 \mcsr/_1272_ ( .A(\mcsr/_0441_ ), .ZN(\mcsr/_0442_ ) );
BUF_X4 \mcsr/_1273_ ( .A(\mcsr/_0376_ ), .Z(\mcsr/_0443_ ) );
OAI21_X1 \mcsr/_1274_ ( .A(\mcsr/_0442_ ), .B1(\mcsr/_0159_ ), .B2(\mcsr/_0443_ ), .ZN(\mcsr/_0444_ ) );
OR2_X1 \mcsr/_1275_ ( .A1(\mcsr/_0421_ ), .A2(\mcsr/_0255_ ), .ZN(\mcsr/_0445_ ) );
INV_X1 \mcsr/_1276_ ( .A(\mcsr/_0223_ ), .ZN(\mcsr/_0446_ ) );
AOI22_X2 \mcsr/_1277_ ( .A1(\mcsr/_0388_ ), .A2(\mcsr/_0446_ ), .B1(\mcsr/_0391_ ), .B2(\mcsr/_0393_ ), .ZN(\mcsr/_0447_ ) );
NAND2_X1 \mcsr/_1278_ ( .A1(\mcsr/_0445_ ), .A2(\mcsr/_0447_ ), .ZN(\mcsr/_0448_ ) );
AOI21_X1 \mcsr/_1279_ ( .A(\mcsr/_0364_ ), .B1(\mcsr/_0444_ ), .B2(\mcsr/_0448_ ), .ZN(\mcsr/_0833_ ) );
OAI211_X2 \mcsr/_1280_ ( .A(\mcsr/_0402_ ), .B(\mcsr/_0403_ ), .C1(\mcsr/_0161_ ), .C2(\mcsr/_0440_ ), .ZN(\mcsr/_0449_ ) );
INV_X1 \mcsr/_1281_ ( .A(\mcsr/_0449_ ), .ZN(\mcsr/_0450_ ) );
OAI21_X1 \mcsr/_1282_ ( .A(\mcsr/_0450_ ), .B1(\mcsr/_0129_ ), .B2(\mcsr/_0443_ ), .ZN(\mcsr/_0451_ ) );
OR2_X1 \mcsr/_1283_ ( .A1(\mcsr/_0421_ ), .A2(\mcsr/_0225_ ), .ZN(\mcsr/_0452_ ) );
INV_X1 \mcsr/_1284_ ( .A(\mcsr/_0193_ ), .ZN(\mcsr/_0453_ ) );
AOI22_X2 \mcsr/_1285_ ( .A1(\mcsr/_0388_ ), .A2(\mcsr/_0453_ ), .B1(\mcsr/_0391_ ), .B2(\mcsr/_0393_ ), .ZN(\mcsr/_0454_ ) );
NAND2_X1 \mcsr/_1286_ ( .A1(\mcsr/_0452_ ), .A2(\mcsr/_0454_ ), .ZN(\mcsr/_0455_ ) );
AOI21_X1 \mcsr/_1287_ ( .A(\mcsr/_0364_ ), .B1(\mcsr/_0451_ ), .B2(\mcsr/_0455_ ), .ZN(\mcsr/_0803_ ) );
OR2_X1 \mcsr/_1288_ ( .A1(\mcsr/_0375_ ), .A2(\mcsr/_0226_ ), .ZN(\mcsr/_0456_ ) );
NOR2_X1 \mcsr/_1289_ ( .A1(\mcsr/_0261_ ), .A2(\mcsr/_0260_ ), .ZN(\mcsr/_0457_ ) );
AND3_X1 \mcsr/_1290_ ( .A1(\mcsr/_0457_ ), .A2(\mcsr/_0340_ ), .A3(\mcsr/_0256_ ), .ZN(\mcsr/_0458_ ) );
NAND3_X1 \mcsr/_1291_ ( .A1(\mcsr/_0355_ ), .A2(\mcsr/_0336_ ), .A3(\mcsr/_0458_ ), .ZN(\mcsr/_0459_ ) );
NAND2_X1 \mcsr/_1292_ ( .A1(\mcsr/_0358_ ), .A2(\mcsr/_0459_ ), .ZN(\mcsr/_0460_ ) );
INV_X1 \mcsr/_1293_ ( .A(\mcsr/_0362_ ), .ZN(\mcsr/_0461_ ) );
OAI211_X2 \mcsr/_1294_ ( .A(\mcsr/_0456_ ), .B(\mcsr/_0460_ ), .C1(\mcsr/_0194_ ), .C2(\mcsr/_0461_ ), .ZN(\mcsr/_0462_ ) );
BUF_X4 \mcsr/_1295_ ( .A(\mcsr/_0352_ ), .Z(\mcsr/_0463_ ) );
INV_X1 \mcsr/_1296_ ( .A(\mcsr/_0463_ ), .ZN(\mcsr/_0464_ ) );
INV_X1 \mcsr/_1297_ ( .A(\mcsr/_0162_ ), .ZN(\mcsr/_0465_ ) );
OAI21_X1 \mcsr/_1298_ ( .A(\mcsr/_0465_ ), .B1(\mcsr/_0342_ ), .B2(\mcsr/_0369_ ), .ZN(\mcsr/_0466_ ) );
OAI211_X2 \mcsr/_1299_ ( .A(\mcsr/_0346_ ), .B(\mcsr/_0466_ ), .C1(\mcsr/_0377_ ), .C2(\mcsr/_0130_ ), .ZN(\mcsr/_0467_ ) );
NAND3_X1 \mcsr/_1300_ ( .A1(\mcsr/_0462_ ), .A2(\mcsr/_0464_ ), .A3(\mcsr/_0467_ ), .ZN(\mcsr/_0804_ ) );
OR2_X1 \mcsr/_1301_ ( .A1(\mcsr/_0375_ ), .A2(\mcsr/_0227_ ), .ZN(\mcsr/_0468_ ) );
OAI211_X2 \mcsr/_1302_ ( .A(\mcsr/_0468_ ), .B(\mcsr/_0460_ ), .C1(\mcsr/_0195_ ), .C2(\mcsr/_0461_ ), .ZN(\mcsr/_0469_ ) );
INV_X1 \mcsr/_1303_ ( .A(\mcsr/_0163_ ), .ZN(\mcsr/_0470_ ) );
OAI21_X1 \mcsr/_1304_ ( .A(\mcsr/_0470_ ), .B1(\mcsr/_0342_ ), .B2(\mcsr/_0369_ ), .ZN(\mcsr/_0471_ ) );
OAI211_X2 \mcsr/_1305_ ( .A(\mcsr/_0346_ ), .B(\mcsr/_0471_ ), .C1(\mcsr/_0377_ ), .C2(\mcsr/_0131_ ), .ZN(\mcsr/_0472_ ) );
NAND3_X1 \mcsr/_1306_ ( .A1(\mcsr/_0469_ ), .A2(\mcsr/_0464_ ), .A3(\mcsr/_0472_ ), .ZN(\mcsr/_0805_ ) );
BUF_X4 \mcsr/_1307_ ( .A(\mcsr/_0352_ ), .Z(\mcsr/_0473_ ) );
OAI211_X2 \mcsr/_1308_ ( .A(\mcsr/_0402_ ), .B(\mcsr/_0403_ ), .C1(\mcsr/_0164_ ), .C2(\mcsr/_0440_ ), .ZN(\mcsr/_0474_ ) );
INV_X1 \mcsr/_1309_ ( .A(\mcsr/_0474_ ), .ZN(\mcsr/_0475_ ) );
OAI21_X1 \mcsr/_1310_ ( .A(\mcsr/_0475_ ), .B1(\mcsr/_0132_ ), .B2(\mcsr/_0443_ ), .ZN(\mcsr/_0476_ ) );
OR2_X1 \mcsr/_1311_ ( .A1(\mcsr/_0421_ ), .A2(\mcsr/_0228_ ), .ZN(\mcsr/_0477_ ) );
INV_X1 \mcsr/_1312_ ( .A(\mcsr/_0196_ ), .ZN(\mcsr/_0478_ ) );
AOI22_X2 \mcsr/_1313_ ( .A1(\mcsr/_0388_ ), .A2(\mcsr/_0478_ ), .B1(\mcsr/_0391_ ), .B2(\mcsr/_0393_ ), .ZN(\mcsr/_0479_ ) );
NAND2_X1 \mcsr/_1314_ ( .A1(\mcsr/_0477_ ), .A2(\mcsr/_0479_ ), .ZN(\mcsr/_0480_ ) );
AOI21_X1 \mcsr/_1315_ ( .A(\mcsr/_0473_ ), .B1(\mcsr/_0476_ ), .B2(\mcsr/_0480_ ), .ZN(\mcsr/_0806_ ) );
OAI211_X2 \mcsr/_1316_ ( .A(\mcsr/_0402_ ), .B(\mcsr/_0403_ ), .C1(\mcsr/_0165_ ), .C2(\mcsr/_0440_ ), .ZN(\mcsr/_0481_ ) );
INV_X1 \mcsr/_1317_ ( .A(\mcsr/_0481_ ), .ZN(\mcsr/_0482_ ) );
OAI21_X1 \mcsr/_1318_ ( .A(\mcsr/_0482_ ), .B1(\mcsr/_0133_ ), .B2(\mcsr/_0443_ ), .ZN(\mcsr/_0483_ ) );
OR2_X1 \mcsr/_1319_ ( .A1(\mcsr/_0421_ ), .A2(\mcsr/_0229_ ), .ZN(\mcsr/_0484_ ) );
INV_X1 \mcsr/_1320_ ( .A(\mcsr/_0197_ ), .ZN(\mcsr/_0485_ ) );
AOI22_X2 \mcsr/_1321_ ( .A1(\mcsr/_0388_ ), .A2(\mcsr/_0485_ ), .B1(\mcsr/_0391_ ), .B2(\mcsr/_0393_ ), .ZN(\mcsr/_0486_ ) );
NAND2_X1 \mcsr/_1322_ ( .A1(\mcsr/_0484_ ), .A2(\mcsr/_0486_ ), .ZN(\mcsr/_0487_ ) );
AOI21_X1 \mcsr/_1323_ ( .A(\mcsr/_0473_ ), .B1(\mcsr/_0483_ ), .B2(\mcsr/_0487_ ), .ZN(\mcsr/_0807_ ) );
OAI211_X2 \mcsr/_1324_ ( .A(\mcsr/_0402_ ), .B(\mcsr/_0403_ ), .C1(\mcsr/_0166_ ), .C2(\mcsr/_0440_ ), .ZN(\mcsr/_0488_ ) );
INV_X1 \mcsr/_1325_ ( .A(\mcsr/_0488_ ), .ZN(\mcsr/_0489_ ) );
OAI21_X1 \mcsr/_1326_ ( .A(\mcsr/_0489_ ), .B1(\mcsr/_0134_ ), .B2(\mcsr/_0443_ ), .ZN(\mcsr/_0490_ ) );
OR2_X1 \mcsr/_1327_ ( .A1(\mcsr/_0421_ ), .A2(\mcsr/_0230_ ), .ZN(\mcsr/_0491_ ) );
BUF_X4 \mcsr/_1328_ ( .A(\mcsr/_0375_ ), .Z(\mcsr/_0492_ ) );
INV_X1 \mcsr/_1329_ ( .A(\mcsr/_0198_ ), .ZN(\mcsr/_0493_ ) );
BUF_X32 \mcsr/_1330_ ( .A(\mcsr/_0390_ ), .Z(\mcsr/_0494_ ) );
BUF_X16 \mcsr/_1331_ ( .A(\mcsr/_0392_ ), .Z(\mcsr/_0495_ ) );
AOI22_X2 \mcsr/_1332_ ( .A1(\mcsr/_0492_ ), .A2(\mcsr/_0493_ ), .B1(\mcsr/_0494_ ), .B2(\mcsr/_0495_ ), .ZN(\mcsr/_0496_ ) );
NAND2_X1 \mcsr/_1333_ ( .A1(\mcsr/_0491_ ), .A2(\mcsr/_0496_ ), .ZN(\mcsr/_0497_ ) );
AOI21_X1 \mcsr/_1334_ ( .A(\mcsr/_0473_ ), .B1(\mcsr/_0490_ ), .B2(\mcsr/_0497_ ), .ZN(\mcsr/_0808_ ) );
BUF_X8 \mcsr/_1335_ ( .A(\mcsr/_0390_ ), .Z(\mcsr/_0498_ ) );
BUF_X8 \mcsr/_1336_ ( .A(\mcsr/_0392_ ), .Z(\mcsr/_0499_ ) );
OAI211_X2 \mcsr/_1337_ ( .A(\mcsr/_0498_ ), .B(\mcsr/_0499_ ), .C1(\mcsr/_0167_ ), .C2(\mcsr/_0440_ ), .ZN(\mcsr/_0500_ ) );
INV_X1 \mcsr/_1338_ ( .A(\mcsr/_0500_ ), .ZN(\mcsr/_0501_ ) );
OAI21_X1 \mcsr/_1339_ ( .A(\mcsr/_0501_ ), .B1(\mcsr/_0135_ ), .B2(\mcsr/_0443_ ), .ZN(\mcsr/_0502_ ) );
OR2_X1 \mcsr/_1340_ ( .A1(\mcsr/_0421_ ), .A2(\mcsr/_0231_ ), .ZN(\mcsr/_0503_ ) );
INV_X1 \mcsr/_1341_ ( .A(\mcsr/_0199_ ), .ZN(\mcsr/_0504_ ) );
AOI22_X2 \mcsr/_1342_ ( .A1(\mcsr/_0492_ ), .A2(\mcsr/_0504_ ), .B1(\mcsr/_0494_ ), .B2(\mcsr/_0495_ ), .ZN(\mcsr/_0505_ ) );
NAND2_X1 \mcsr/_1343_ ( .A1(\mcsr/_0503_ ), .A2(\mcsr/_0505_ ), .ZN(\mcsr/_0506_ ) );
AOI21_X1 \mcsr/_1344_ ( .A(\mcsr/_0473_ ), .B1(\mcsr/_0502_ ), .B2(\mcsr/_0506_ ), .ZN(\mcsr/_0809_ ) );
OAI211_X2 \mcsr/_1345_ ( .A(\mcsr/_0498_ ), .B(\mcsr/_0499_ ), .C1(\mcsr/_0168_ ), .C2(\mcsr/_0440_ ), .ZN(\mcsr/_0507_ ) );
INV_X1 \mcsr/_1346_ ( .A(\mcsr/_0507_ ), .ZN(\mcsr/_0508_ ) );
OAI21_X1 \mcsr/_1347_ ( .A(\mcsr/_0508_ ), .B1(\mcsr/_0136_ ), .B2(\mcsr/_0443_ ), .ZN(\mcsr/_0509_ ) );
OR2_X1 \mcsr/_1348_ ( .A1(\mcsr/_0421_ ), .A2(\mcsr/_0232_ ), .ZN(\mcsr/_0510_ ) );
INV_X1 \mcsr/_1349_ ( .A(\mcsr/_0200_ ), .ZN(\mcsr/_0511_ ) );
AOI22_X2 \mcsr/_1350_ ( .A1(\mcsr/_0492_ ), .A2(\mcsr/_0511_ ), .B1(\mcsr/_0494_ ), .B2(\mcsr/_0495_ ), .ZN(\mcsr/_0512_ ) );
NAND2_X1 \mcsr/_1351_ ( .A1(\mcsr/_0510_ ), .A2(\mcsr/_0512_ ), .ZN(\mcsr/_0513_ ) );
AOI21_X1 \mcsr/_1352_ ( .A(\mcsr/_0473_ ), .B1(\mcsr/_0509_ ), .B2(\mcsr/_0513_ ), .ZN(\mcsr/_0810_ ) );
OAI211_X2 \mcsr/_1353_ ( .A(\mcsr/_0498_ ), .B(\mcsr/_0499_ ), .C1(\mcsr/_0169_ ), .C2(\mcsr/_0440_ ), .ZN(\mcsr/_0514_ ) );
INV_X1 \mcsr/_1354_ ( .A(\mcsr/_0514_ ), .ZN(\mcsr/_0515_ ) );
OAI21_X1 \mcsr/_1355_ ( .A(\mcsr/_0515_ ), .B1(\mcsr/_0137_ ), .B2(\mcsr/_0443_ ), .ZN(\mcsr/_0516_ ) );
CLKBUF_X2 \mcsr/_1356_ ( .A(\mcsr/_0374_ ), .Z(\mcsr/_0517_ ) );
OR2_X1 \mcsr/_1357_ ( .A1(\mcsr/_0517_ ), .A2(\mcsr/_0233_ ), .ZN(\mcsr/_0518_ ) );
INV_X1 \mcsr/_1358_ ( .A(\mcsr/_0201_ ), .ZN(\mcsr/_0519_ ) );
AOI22_X2 \mcsr/_1359_ ( .A1(\mcsr/_0492_ ), .A2(\mcsr/_0519_ ), .B1(\mcsr/_0494_ ), .B2(\mcsr/_0495_ ), .ZN(\mcsr/_0520_ ) );
NAND2_X1 \mcsr/_1360_ ( .A1(\mcsr/_0518_ ), .A2(\mcsr/_0520_ ), .ZN(\mcsr/_0521_ ) );
AOI21_X1 \mcsr/_1361_ ( .A(\mcsr/_0473_ ), .B1(\mcsr/_0516_ ), .B2(\mcsr/_0521_ ), .ZN(\mcsr/_0811_ ) );
OAI211_X2 \mcsr/_1362_ ( .A(\mcsr/_0498_ ), .B(\mcsr/_0499_ ), .C1(\mcsr/_0170_ ), .C2(\mcsr/_0440_ ), .ZN(\mcsr/_0522_ ) );
INV_X1 \mcsr/_1363_ ( .A(\mcsr/_0522_ ), .ZN(\mcsr/_0523_ ) );
OAI21_X1 \mcsr/_1364_ ( .A(\mcsr/_0523_ ), .B1(\mcsr/_0138_ ), .B2(\mcsr/_0443_ ), .ZN(\mcsr/_0524_ ) );
OR2_X1 \mcsr/_1365_ ( .A1(\mcsr/_0517_ ), .A2(\mcsr/_0234_ ), .ZN(\mcsr/_0525_ ) );
INV_X1 \mcsr/_1366_ ( .A(\mcsr/_0202_ ), .ZN(\mcsr/_0526_ ) );
AOI22_X2 \mcsr/_1367_ ( .A1(\mcsr/_0492_ ), .A2(\mcsr/_0526_ ), .B1(\mcsr/_0494_ ), .B2(\mcsr/_0495_ ), .ZN(\mcsr/_0527_ ) );
NAND2_X1 \mcsr/_1368_ ( .A1(\mcsr/_0525_ ), .A2(\mcsr/_0527_ ), .ZN(\mcsr/_0528_ ) );
AOI21_X1 \mcsr/_1369_ ( .A(\mcsr/_0473_ ), .B1(\mcsr/_0524_ ), .B2(\mcsr/_0528_ ), .ZN(\mcsr/_0812_ ) );
OAI211_X2 \mcsr/_1370_ ( .A(\mcsr/_0498_ ), .B(\mcsr/_0499_ ), .C1(\mcsr/_0172_ ), .C2(\mcsr/_0440_ ), .ZN(\mcsr/_0529_ ) );
INV_X1 \mcsr/_1371_ ( .A(\mcsr/_0529_ ), .ZN(\mcsr/_0530_ ) );
OAI21_X1 \mcsr/_1372_ ( .A(\mcsr/_0530_ ), .B1(\mcsr/_0140_ ), .B2(\mcsr/_0443_ ), .ZN(\mcsr/_0531_ ) );
OR2_X1 \mcsr/_1373_ ( .A1(\mcsr/_0517_ ), .A2(\mcsr/_0236_ ), .ZN(\mcsr/_0532_ ) );
INV_X1 \mcsr/_1374_ ( .A(\mcsr/_0204_ ), .ZN(\mcsr/_0533_ ) );
AOI22_X2 \mcsr/_1375_ ( .A1(\mcsr/_0492_ ), .A2(\mcsr/_0533_ ), .B1(\mcsr/_0494_ ), .B2(\mcsr/_0495_ ), .ZN(\mcsr/_0534_ ) );
NAND2_X1 \mcsr/_1376_ ( .A1(\mcsr/_0532_ ), .A2(\mcsr/_0534_ ), .ZN(\mcsr/_0535_ ) );
AOI21_X1 \mcsr/_1377_ ( .A(\mcsr/_0473_ ), .B1(\mcsr/_0531_ ), .B2(\mcsr/_0535_ ), .ZN(\mcsr/_0814_ ) );
BUF_X8 \mcsr/_1378_ ( .A(\mcsr/_0370_ ), .Z(\mcsr/_0536_ ) );
OAI211_X2 \mcsr/_1379_ ( .A(\mcsr/_0498_ ), .B(\mcsr/_0499_ ), .C1(\mcsr/_0173_ ), .C2(\mcsr/_0536_ ), .ZN(\mcsr/_0537_ ) );
INV_X1 \mcsr/_1380_ ( .A(\mcsr/_0537_ ), .ZN(\mcsr/_0538_ ) );
BUF_X4 \mcsr/_1381_ ( .A(\mcsr/_0376_ ), .Z(\mcsr/_0539_ ) );
OAI21_X1 \mcsr/_1382_ ( .A(\mcsr/_0538_ ), .B1(\mcsr/_0141_ ), .B2(\mcsr/_0539_ ), .ZN(\mcsr/_0540_ ) );
OR2_X1 \mcsr/_1383_ ( .A1(\mcsr/_0517_ ), .A2(\mcsr/_0237_ ), .ZN(\mcsr/_0541_ ) );
INV_X1 \mcsr/_1384_ ( .A(\mcsr/_0205_ ), .ZN(\mcsr/_0542_ ) );
AOI22_X2 \mcsr/_1385_ ( .A1(\mcsr/_0492_ ), .A2(\mcsr/_0542_ ), .B1(\mcsr/_0494_ ), .B2(\mcsr/_0495_ ), .ZN(\mcsr/_0543_ ) );
NAND2_X1 \mcsr/_1386_ ( .A1(\mcsr/_0541_ ), .A2(\mcsr/_0543_ ), .ZN(\mcsr/_0544_ ) );
AOI21_X1 \mcsr/_1387_ ( .A(\mcsr/_0473_ ), .B1(\mcsr/_0540_ ), .B2(\mcsr/_0544_ ), .ZN(\mcsr/_0815_ ) );
OAI211_X2 \mcsr/_1388_ ( .A(\mcsr/_0498_ ), .B(\mcsr/_0499_ ), .C1(\mcsr/_0174_ ), .C2(\mcsr/_0536_ ), .ZN(\mcsr/_0545_ ) );
INV_X1 \mcsr/_1389_ ( .A(\mcsr/_0545_ ), .ZN(\mcsr/_0546_ ) );
OAI21_X1 \mcsr/_1390_ ( .A(\mcsr/_0546_ ), .B1(\mcsr/_0142_ ), .B2(\mcsr/_0539_ ), .ZN(\mcsr/_0547_ ) );
OR2_X1 \mcsr/_1391_ ( .A1(\mcsr/_0517_ ), .A2(\mcsr/_0238_ ), .ZN(\mcsr/_0548_ ) );
INV_X1 \mcsr/_1392_ ( .A(\mcsr/_0206_ ), .ZN(\mcsr/_0549_ ) );
AOI22_X2 \mcsr/_1393_ ( .A1(\mcsr/_0492_ ), .A2(\mcsr/_0549_ ), .B1(\mcsr/_0494_ ), .B2(\mcsr/_0495_ ), .ZN(\mcsr/_0550_ ) );
NAND2_X1 \mcsr/_1394_ ( .A1(\mcsr/_0548_ ), .A2(\mcsr/_0550_ ), .ZN(\mcsr/_0551_ ) );
AOI21_X1 \mcsr/_1395_ ( .A(\mcsr/_0473_ ), .B1(\mcsr/_0547_ ), .B2(\mcsr/_0551_ ), .ZN(\mcsr/_0816_ ) );
OAI211_X2 \mcsr/_1396_ ( .A(\mcsr/_0498_ ), .B(\mcsr/_0499_ ), .C1(\mcsr/_0175_ ), .C2(\mcsr/_0536_ ), .ZN(\mcsr/_0552_ ) );
INV_X1 \mcsr/_1397_ ( .A(\mcsr/_0552_ ), .ZN(\mcsr/_0553_ ) );
OAI21_X1 \mcsr/_1398_ ( .A(\mcsr/_0553_ ), .B1(\mcsr/_0143_ ), .B2(\mcsr/_0539_ ), .ZN(\mcsr/_0554_ ) );
OR2_X1 \mcsr/_1399_ ( .A1(\mcsr/_0517_ ), .A2(\mcsr/_0239_ ), .ZN(\mcsr/_0555_ ) );
INV_X1 \mcsr/_1400_ ( .A(\mcsr/_0207_ ), .ZN(\mcsr/_0556_ ) );
AOI22_X2 \mcsr/_1401_ ( .A1(\mcsr/_0492_ ), .A2(\mcsr/_0556_ ), .B1(\mcsr/_0494_ ), .B2(\mcsr/_0495_ ), .ZN(\mcsr/_0557_ ) );
NAND2_X1 \mcsr/_1402_ ( .A1(\mcsr/_0555_ ), .A2(\mcsr/_0557_ ), .ZN(\mcsr/_0558_ ) );
AOI21_X1 \mcsr/_1403_ ( .A(\mcsr/_0463_ ), .B1(\mcsr/_0554_ ), .B2(\mcsr/_0558_ ), .ZN(\mcsr/_0817_ ) );
OAI211_X2 \mcsr/_1404_ ( .A(\mcsr/_0498_ ), .B(\mcsr/_0499_ ), .C1(\mcsr/_0176_ ), .C2(\mcsr/_0536_ ), .ZN(\mcsr/_0559_ ) );
INV_X1 \mcsr/_1405_ ( .A(\mcsr/_0559_ ), .ZN(\mcsr/_0560_ ) );
OAI21_X1 \mcsr/_1406_ ( .A(\mcsr/_0560_ ), .B1(\mcsr/_0144_ ), .B2(\mcsr/_0539_ ), .ZN(\mcsr/_0561_ ) );
OR2_X1 \mcsr/_1407_ ( .A1(\mcsr/_0517_ ), .A2(\mcsr/_0240_ ), .ZN(\mcsr/_0562_ ) );
INV_X1 \mcsr/_1408_ ( .A(\mcsr/_0208_ ), .ZN(\mcsr/_0563_ ) );
AOI22_X2 \mcsr/_1409_ ( .A1(\mcsr/_0492_ ), .A2(\mcsr/_0563_ ), .B1(\mcsr/_0494_ ), .B2(\mcsr/_0495_ ), .ZN(\mcsr/_0564_ ) );
NAND2_X1 \mcsr/_1410_ ( .A1(\mcsr/_0562_ ), .A2(\mcsr/_0564_ ), .ZN(\mcsr/_0565_ ) );
AOI21_X1 \mcsr/_1411_ ( .A(\mcsr/_0463_ ), .B1(\mcsr/_0561_ ), .B2(\mcsr/_0565_ ), .ZN(\mcsr/_0818_ ) );
OAI211_X2 \mcsr/_1412_ ( .A(\mcsr/_0498_ ), .B(\mcsr/_0499_ ), .C1(\mcsr/_0177_ ), .C2(\mcsr/_0536_ ), .ZN(\mcsr/_0566_ ) );
INV_X1 \mcsr/_1413_ ( .A(\mcsr/_0566_ ), .ZN(\mcsr/_0567_ ) );
OAI21_X1 \mcsr/_1414_ ( .A(\mcsr/_0567_ ), .B1(\mcsr/_0145_ ), .B2(\mcsr/_0539_ ), .ZN(\mcsr/_0568_ ) );
OR2_X1 \mcsr/_1415_ ( .A1(\mcsr/_0517_ ), .A2(\mcsr/_0241_ ), .ZN(\mcsr/_0569_ ) );
INV_X1 \mcsr/_1416_ ( .A(\mcsr/_0209_ ), .ZN(\mcsr/_0570_ ) );
AOI22_X1 \mcsr/_1417_ ( .A1(\mcsr/_0386_ ), .A2(\mcsr/_0570_ ), .B1(\mcsr/_0366_ ), .B2(\mcsr/_0368_ ), .ZN(\mcsr/_0571_ ) );
NAND2_X1 \mcsr/_1418_ ( .A1(\mcsr/_0569_ ), .A2(\mcsr/_0571_ ), .ZN(\mcsr/_0572_ ) );
AOI21_X1 \mcsr/_1419_ ( .A(\mcsr/_0463_ ), .B1(\mcsr/_0568_ ), .B2(\mcsr/_0572_ ), .ZN(\mcsr/_0819_ ) );
OAI211_X2 \mcsr/_1420_ ( .A(\mcsr/_0390_ ), .B(\mcsr/_0392_ ), .C1(\mcsr/_0178_ ), .C2(\mcsr/_0536_ ), .ZN(\mcsr/_0573_ ) );
INV_X1 \mcsr/_1421_ ( .A(\mcsr/_0573_ ), .ZN(\mcsr/_0574_ ) );
OAI21_X1 \mcsr/_1422_ ( .A(\mcsr/_0574_ ), .B1(\mcsr/_0146_ ), .B2(\mcsr/_0539_ ), .ZN(\mcsr/_0575_ ) );
OR2_X1 \mcsr/_1423_ ( .A1(\mcsr/_0517_ ), .A2(\mcsr/_0242_ ), .ZN(\mcsr/_0576_ ) );
INV_X1 \mcsr/_1424_ ( .A(\mcsr/_0210_ ), .ZN(\mcsr/_0577_ ) );
AOI22_X1 \mcsr/_1425_ ( .A1(\mcsr/_0386_ ), .A2(\mcsr/_0577_ ), .B1(\mcsr/_0366_ ), .B2(\mcsr/_0368_ ), .ZN(\mcsr/_0578_ ) );
NAND2_X1 \mcsr/_1426_ ( .A1(\mcsr/_0576_ ), .A2(\mcsr/_0578_ ), .ZN(\mcsr/_0579_ ) );
AOI21_X1 \mcsr/_1427_ ( .A(\mcsr/_0463_ ), .B1(\mcsr/_0575_ ), .B2(\mcsr/_0579_ ), .ZN(\mcsr/_0820_ ) );
OAI211_X2 \mcsr/_1428_ ( .A(\mcsr/_0390_ ), .B(\mcsr/_0392_ ), .C1(\mcsr/_0179_ ), .C2(\mcsr/_0536_ ), .ZN(\mcsr/_0580_ ) );
INV_X1 \mcsr/_1429_ ( .A(\mcsr/_0580_ ), .ZN(\mcsr/_0581_ ) );
OAI21_X1 \mcsr/_1430_ ( .A(\mcsr/_0581_ ), .B1(\mcsr/_0147_ ), .B2(\mcsr/_0539_ ), .ZN(\mcsr/_0582_ ) );
OR2_X1 \mcsr/_1431_ ( .A1(\mcsr/_0517_ ), .A2(\mcsr/_0243_ ), .ZN(\mcsr/_0583_ ) );
INV_X1 \mcsr/_1432_ ( .A(\mcsr/_0211_ ), .ZN(\mcsr/_0584_ ) );
AOI22_X1 \mcsr/_1433_ ( .A1(\mcsr/_0386_ ), .A2(\mcsr/_0584_ ), .B1(\mcsr/_0366_ ), .B2(\mcsr/_0368_ ), .ZN(\mcsr/_0585_ ) );
NAND2_X1 \mcsr/_1434_ ( .A1(\mcsr/_0583_ ), .A2(\mcsr/_0585_ ), .ZN(\mcsr/_0586_ ) );
AOI21_X1 \mcsr/_1435_ ( .A(\mcsr/_0463_ ), .B1(\mcsr/_0582_ ), .B2(\mcsr/_0586_ ), .ZN(\mcsr/_0821_ ) );
OAI211_X2 \mcsr/_1436_ ( .A(\mcsr/_0390_ ), .B(\mcsr/_0392_ ), .C1(\mcsr/_0180_ ), .C2(\mcsr/_0536_ ), .ZN(\mcsr/_0587_ ) );
INV_X1 \mcsr/_1437_ ( .A(\mcsr/_0587_ ), .ZN(\mcsr/_0588_ ) );
OAI21_X1 \mcsr/_1438_ ( .A(\mcsr/_0588_ ), .B1(\mcsr/_0148_ ), .B2(\mcsr/_0539_ ), .ZN(\mcsr/_0589_ ) );
OR2_X1 \mcsr/_1439_ ( .A1(\mcsr/_0375_ ), .A2(\mcsr/_0244_ ), .ZN(\mcsr/_0590_ ) );
INV_X1 \mcsr/_1440_ ( .A(\mcsr/_0212_ ), .ZN(\mcsr/_0591_ ) );
AOI22_X1 \mcsr/_1441_ ( .A1(\mcsr/_0386_ ), .A2(\mcsr/_0591_ ), .B1(\mcsr/_0366_ ), .B2(\mcsr/_0368_ ), .ZN(\mcsr/_0592_ ) );
NAND2_X1 \mcsr/_1442_ ( .A1(\mcsr/_0590_ ), .A2(\mcsr/_0592_ ), .ZN(\mcsr/_0593_ ) );
AOI21_X1 \mcsr/_1443_ ( .A(\mcsr/_0463_ ), .B1(\mcsr/_0589_ ), .B2(\mcsr/_0593_ ), .ZN(\mcsr/_0822_ ) );
OAI211_X2 \mcsr/_1444_ ( .A(\mcsr/_0390_ ), .B(\mcsr/_0392_ ), .C1(\mcsr/_0181_ ), .C2(\mcsr/_0536_ ), .ZN(\mcsr/_0594_ ) );
INV_X1 \mcsr/_1445_ ( .A(\mcsr/_0594_ ), .ZN(\mcsr/_0595_ ) );
OAI21_X1 \mcsr/_1446_ ( .A(\mcsr/_0595_ ), .B1(\mcsr/_0149_ ), .B2(\mcsr/_0539_ ), .ZN(\mcsr/_0596_ ) );
OR2_X1 \mcsr/_1447_ ( .A1(\mcsr/_0375_ ), .A2(\mcsr/_0245_ ), .ZN(\mcsr/_0597_ ) );
INV_X1 \mcsr/_1448_ ( .A(\mcsr/_0213_ ), .ZN(\mcsr/_0598_ ) );
AOI22_X1 \mcsr/_1449_ ( .A1(\mcsr/_0386_ ), .A2(\mcsr/_0598_ ), .B1(\mcsr/_0366_ ), .B2(\mcsr/_0368_ ), .ZN(\mcsr/_0599_ ) );
NAND2_X1 \mcsr/_1450_ ( .A1(\mcsr/_0597_ ), .A2(\mcsr/_0599_ ), .ZN(\mcsr/_0600_ ) );
AOI21_X1 \mcsr/_1451_ ( .A(\mcsr/_0463_ ), .B1(\mcsr/_0596_ ), .B2(\mcsr/_0600_ ), .ZN(\mcsr/_0823_ ) );
OAI211_X2 \mcsr/_1452_ ( .A(\mcsr/_0390_ ), .B(\mcsr/_0392_ ), .C1(\mcsr/_0183_ ), .C2(\mcsr/_0536_ ), .ZN(\mcsr/_0601_ ) );
INV_X1 \mcsr/_1453_ ( .A(\mcsr/_0601_ ), .ZN(\mcsr/_0602_ ) );
OAI21_X1 \mcsr/_1454_ ( .A(\mcsr/_0602_ ), .B1(\mcsr/_0151_ ), .B2(\mcsr/_0539_ ), .ZN(\mcsr/_0603_ ) );
OR2_X1 \mcsr/_1455_ ( .A1(\mcsr/_0375_ ), .A2(\mcsr/_0247_ ), .ZN(\mcsr/_0604_ ) );
INV_X1 \mcsr/_1456_ ( .A(\mcsr/_0215_ ), .ZN(\mcsr/_0605_ ) );
AOI22_X1 \mcsr/_1457_ ( .A1(\mcsr/_0386_ ), .A2(\mcsr/_0605_ ), .B1(\mcsr/_0366_ ), .B2(\mcsr/_0368_ ), .ZN(\mcsr/_0606_ ) );
NAND2_X1 \mcsr/_1458_ ( .A1(\mcsr/_0604_ ), .A2(\mcsr/_0606_ ), .ZN(\mcsr/_0607_ ) );
AOI21_X1 \mcsr/_1459_ ( .A(\mcsr/_0463_ ), .B1(\mcsr/_0603_ ), .B2(\mcsr/_0607_ ), .ZN(\mcsr/_0825_ ) );
OAI211_X2 \mcsr/_1460_ ( .A(\mcsr/_0390_ ), .B(\mcsr/_0392_ ), .C1(\mcsr/_0184_ ), .C2(\mcsr/_0370_ ), .ZN(\mcsr/_0608_ ) );
INV_X1 \mcsr/_1461_ ( .A(\mcsr/_0608_ ), .ZN(\mcsr/_0609_ ) );
OAI21_X1 \mcsr/_1462_ ( .A(\mcsr/_0609_ ), .B1(\mcsr/_0152_ ), .B2(\mcsr/_0376_ ), .ZN(\mcsr/_0610_ ) );
OR2_X1 \mcsr/_1463_ ( .A1(\mcsr/_0375_ ), .A2(\mcsr/_0248_ ), .ZN(\mcsr/_0611_ ) );
INV_X1 \mcsr/_1464_ ( .A(\mcsr/_0216_ ), .ZN(\mcsr/_0612_ ) );
AOI22_X1 \mcsr/_1465_ ( .A1(\mcsr/_0386_ ), .A2(\mcsr/_0612_ ), .B1(\mcsr/_0366_ ), .B2(\mcsr/_0368_ ), .ZN(\mcsr/_0613_ ) );
NAND2_X1 \mcsr/_1466_ ( .A1(\mcsr/_0611_ ), .A2(\mcsr/_0613_ ), .ZN(\mcsr/_0614_ ) );
AOI21_X1 \mcsr/_1467_ ( .A(\mcsr/_0463_ ), .B1(\mcsr/_0610_ ), .B2(\mcsr/_0614_ ), .ZN(\mcsr/_0826_ ) );
INV_X4 \mcsr/_1468_ ( .A(\mcsr/_0269_ ), .ZN(\mcsr/_0615_ ) );
INV_X2 \mcsr/_1469_ ( .A(\mcsr/_0270_ ), .ZN(\mcsr/_0616_ ) );
BUF_X4 \mcsr/_1470_ ( .A(\mcsr/_0616_ ), .Z(\mcsr/_0617_ ) );
NAND4_X1 \mcsr/_1471_ ( .A1(\mcsr/_0615_ ), .A2(\mcsr/_0617_ ), .A3(\mcsr/_0268_ ), .A4(\mcsr/_0192_ ), .ZN(\mcsr/_0618_ ) );
INV_X32 \mcsr/_1472_ ( .A(\mcsr/_0268_ ), .ZN(\mcsr/_0619_ ) );
BUF_X4 \mcsr/_1473_ ( .A(\mcsr/_0619_ ), .Z(\mcsr/_0620_ ) );
NAND4_X1 \mcsr/_1474_ ( .A1(\mcsr/_0620_ ), .A2(\mcsr/_0617_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0160_ ), .ZN(\mcsr/_0621_ ) );
NAND2_X1 \mcsr/_1475_ ( .A1(\mcsr/_0618_ ), .A2(\mcsr/_0621_ ), .ZN(\mcsr/_0834_ ) );
NAND4_X1 \mcsr/_1476_ ( .A1(\mcsr/_0620_ ), .A2(\mcsr/_0617_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0171_ ), .ZN(\mcsr/_0622_ ) );
NAND4_X1 \mcsr/_1477_ ( .A1(\mcsr/_0615_ ), .A2(\mcsr/_0617_ ), .A3(\mcsr/_0268_ ), .A4(\mcsr/_0203_ ), .ZN(\mcsr/_0623_ ) );
NAND2_X1 \mcsr/_1478_ ( .A1(\mcsr/_0622_ ), .A2(\mcsr/_0623_ ), .ZN(\mcsr/_0845_ ) );
NAND4_X1 \mcsr/_1479_ ( .A1(\mcsr/_0620_ ), .A2(\mcsr/_0617_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0182_ ), .ZN(\mcsr/_0624_ ) );
NOR2_X1 \mcsr/_1480_ ( .A1(\mcsr/_0619_ ), .A2(\mcsr/_0270_ ), .ZN(\mcsr/_0625_ ) );
NAND2_X2 \mcsr/_1481_ ( .A1(\mcsr/_0625_ ), .A2(\mcsr/_0615_ ), .ZN(\mcsr/_0626_ ) );
BUF_X4 \mcsr/_1482_ ( .A(\mcsr/_0626_ ), .Z(\mcsr/_0627_ ) );
OAI21_X1 \mcsr/_1483_ ( .A(\mcsr/_0624_ ), .B1(\mcsr/_0627_ ), .B2(\mcsr/_0389_ ), .ZN(\mcsr/_0856_ ) );
NAND4_X1 \mcsr/_1484_ ( .A1(\mcsr/_0620_ ), .A2(\mcsr/_0617_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0185_ ), .ZN(\mcsr/_0628_ ) );
NAND4_X1 \mcsr/_1485_ ( .A1(\mcsr/_0615_ ), .A2(\mcsr/_0617_ ), .A3(\mcsr/_0268_ ), .A4(\mcsr/_0217_ ), .ZN(\mcsr/_0629_ ) );
NAND2_X1 \mcsr/_1486_ ( .A1(\mcsr/_0628_ ), .A2(\mcsr/_0629_ ), .ZN(\mcsr/_0859_ ) );
NAND4_X1 \mcsr/_1487_ ( .A1(\mcsr/_0620_ ), .A2(\mcsr/_0617_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0186_ ), .ZN(\mcsr/_0630_ ) );
OAI21_X1 \mcsr/_1488_ ( .A(\mcsr/_0630_ ), .B1(\mcsr/_0627_ ), .B2(\mcsr/_0408_ ), .ZN(\mcsr/_0860_ ) );
NAND4_X1 \mcsr/_1489_ ( .A1(\mcsr/_0620_ ), .A2(\mcsr/_0617_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0187_ ), .ZN(\mcsr/_0631_ ) );
OAI21_X1 \mcsr/_1490_ ( .A(\mcsr/_0631_ ), .B1(\mcsr/_0627_ ), .B2(\mcsr/_0415_ ), .ZN(\mcsr/_0861_ ) );
NAND4_X1 \mcsr/_1491_ ( .A1(\mcsr/_0620_ ), .A2(\mcsr/_0617_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0188_ ), .ZN(\mcsr/_0632_ ) );
OAI21_X1 \mcsr/_1492_ ( .A(\mcsr/_0632_ ), .B1(\mcsr/_0627_ ), .B2(\mcsr/_0423_ ), .ZN(\mcsr/_0862_ ) );
BUF_X4 \mcsr/_1493_ ( .A(\mcsr/_0616_ ), .Z(\mcsr/_0633_ ) );
NAND4_X1 \mcsr/_1494_ ( .A1(\mcsr/_0620_ ), .A2(\mcsr/_0633_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0189_ ), .ZN(\mcsr/_0634_ ) );
OAI21_X1 \mcsr/_1495_ ( .A(\mcsr/_0634_ ), .B1(\mcsr/_0627_ ), .B2(\mcsr/_0430_ ), .ZN(\mcsr/_0863_ ) );
NAND4_X1 \mcsr/_1496_ ( .A1(\mcsr/_0620_ ), .A2(\mcsr/_0633_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0190_ ), .ZN(\mcsr/_0635_ ) );
OAI21_X1 \mcsr/_1497_ ( .A(\mcsr/_0635_ ), .B1(\mcsr/_0627_ ), .B2(\mcsr/_0437_ ), .ZN(\mcsr/_0864_ ) );
BUF_X4 \mcsr/_1498_ ( .A(\mcsr/_0619_ ), .Z(\mcsr/_0636_ ) );
NAND4_X1 \mcsr/_1499_ ( .A1(\mcsr/_0636_ ), .A2(\mcsr/_0633_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0191_ ), .ZN(\mcsr/_0637_ ) );
OAI21_X1 \mcsr/_1500_ ( .A(\mcsr/_0637_ ), .B1(\mcsr/_0627_ ), .B2(\mcsr/_0446_ ), .ZN(\mcsr/_0865_ ) );
NAND4_X1 \mcsr/_1501_ ( .A1(\mcsr/_0636_ ), .A2(\mcsr/_0633_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0161_ ), .ZN(\mcsr/_0638_ ) );
OAI21_X1 \mcsr/_1502_ ( .A(\mcsr/_0638_ ), .B1(\mcsr/_0627_ ), .B2(\mcsr/_0453_ ), .ZN(\mcsr/_0835_ ) );
NAND4_X1 \mcsr/_1503_ ( .A1(\mcsr/_0615_ ), .A2(\mcsr/_0633_ ), .A3(\mcsr/_0268_ ), .A4(\mcsr/_0194_ ), .ZN(\mcsr/_0639_ ) );
NOR2_X1 \mcsr/_1504_ ( .A1(\mcsr/_0615_ ), .A2(\mcsr/_0270_ ), .ZN(\mcsr/_0640_ ) );
BUF_X4 \mcsr/_1505_ ( .A(\mcsr/_0640_ ), .Z(\mcsr/_0641_ ) );
NAND2_X1 \mcsr/_1506_ ( .A1(\mcsr/_0641_ ), .A2(\mcsr/_0620_ ), .ZN(\mcsr/_0642_ ) );
OAI21_X1 \mcsr/_1507_ ( .A(\mcsr/_0639_ ), .B1(\mcsr/_0642_ ), .B2(\mcsr/_0465_ ), .ZN(\mcsr/_0836_ ) );
NAND4_X1 \mcsr/_1508_ ( .A1(\mcsr/_0615_ ), .A2(\mcsr/_0633_ ), .A3(\mcsr/_0268_ ), .A4(\mcsr/_0195_ ), .ZN(\mcsr/_0643_ ) );
OAI21_X1 \mcsr/_1509_ ( .A(\mcsr/_0643_ ), .B1(\mcsr/_0642_ ), .B2(\mcsr/_0470_ ), .ZN(\mcsr/_0837_ ) );
NAND4_X1 \mcsr/_1510_ ( .A1(\mcsr/_0636_ ), .A2(\mcsr/_0633_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0164_ ), .ZN(\mcsr/_0644_ ) );
OAI21_X1 \mcsr/_1511_ ( .A(\mcsr/_0644_ ), .B1(\mcsr/_0627_ ), .B2(\mcsr/_0478_ ), .ZN(\mcsr/_0838_ ) );
NAND4_X1 \mcsr/_1512_ ( .A1(\mcsr/_0636_ ), .A2(\mcsr/_0633_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0165_ ), .ZN(\mcsr/_0645_ ) );
OAI21_X1 \mcsr/_1513_ ( .A(\mcsr/_0645_ ), .B1(\mcsr/_0627_ ), .B2(\mcsr/_0485_ ), .ZN(\mcsr/_0839_ ) );
NAND4_X1 \mcsr/_1514_ ( .A1(\mcsr/_0636_ ), .A2(\mcsr/_0633_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0166_ ), .ZN(\mcsr/_0646_ ) );
BUF_X4 \mcsr/_1515_ ( .A(\mcsr/_0626_ ), .Z(\mcsr/_0647_ ) );
OAI21_X1 \mcsr/_1516_ ( .A(\mcsr/_0646_ ), .B1(\mcsr/_0647_ ), .B2(\mcsr/_0493_ ), .ZN(\mcsr/_0840_ ) );
NAND4_X1 \mcsr/_1517_ ( .A1(\mcsr/_0636_ ), .A2(\mcsr/_0633_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0167_ ), .ZN(\mcsr/_0648_ ) );
OAI21_X1 \mcsr/_1518_ ( .A(\mcsr/_0648_ ), .B1(\mcsr/_0647_ ), .B2(\mcsr/_0504_ ), .ZN(\mcsr/_0841_ ) );
BUF_X4 \mcsr/_1519_ ( .A(\mcsr/_0616_ ), .Z(\mcsr/_0649_ ) );
NAND4_X1 \mcsr/_1520_ ( .A1(\mcsr/_0636_ ), .A2(\mcsr/_0649_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0168_ ), .ZN(\mcsr/_0650_ ) );
OAI21_X1 \mcsr/_1521_ ( .A(\mcsr/_0650_ ), .B1(\mcsr/_0647_ ), .B2(\mcsr/_0511_ ), .ZN(\mcsr/_0842_ ) );
NAND4_X1 \mcsr/_1522_ ( .A1(\mcsr/_0636_ ), .A2(\mcsr/_0649_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0169_ ), .ZN(\mcsr/_0651_ ) );
OAI21_X1 \mcsr/_1523_ ( .A(\mcsr/_0651_ ), .B1(\mcsr/_0647_ ), .B2(\mcsr/_0519_ ), .ZN(\mcsr/_0843_ ) );
NAND4_X1 \mcsr/_1524_ ( .A1(\mcsr/_0636_ ), .A2(\mcsr/_0649_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0170_ ), .ZN(\mcsr/_0652_ ) );
OAI21_X1 \mcsr/_1525_ ( .A(\mcsr/_0652_ ), .B1(\mcsr/_0647_ ), .B2(\mcsr/_0526_ ), .ZN(\mcsr/_0844_ ) );
NAND4_X1 \mcsr/_1526_ ( .A1(\mcsr/_0636_ ), .A2(\mcsr/_0649_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0172_ ), .ZN(\mcsr/_0653_ ) );
OAI21_X1 \mcsr/_1527_ ( .A(\mcsr/_0653_ ), .B1(\mcsr/_0647_ ), .B2(\mcsr/_0533_ ), .ZN(\mcsr/_0846_ ) );
BUF_X4 \mcsr/_1528_ ( .A(\mcsr/_0619_ ), .Z(\mcsr/_0654_ ) );
NAND4_X1 \mcsr/_1529_ ( .A1(\mcsr/_0654_ ), .A2(\mcsr/_0649_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0173_ ), .ZN(\mcsr/_0655_ ) );
OAI21_X1 \mcsr/_1530_ ( .A(\mcsr/_0655_ ), .B1(\mcsr/_0647_ ), .B2(\mcsr/_0542_ ), .ZN(\mcsr/_0847_ ) );
NAND4_X1 \mcsr/_1531_ ( .A1(\mcsr/_0654_ ), .A2(\mcsr/_0649_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0174_ ), .ZN(\mcsr/_0656_ ) );
OAI21_X1 \mcsr/_1532_ ( .A(\mcsr/_0656_ ), .B1(\mcsr/_0647_ ), .B2(\mcsr/_0549_ ), .ZN(\mcsr/_0848_ ) );
NAND4_X1 \mcsr/_1533_ ( .A1(\mcsr/_0654_ ), .A2(\mcsr/_0649_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0175_ ), .ZN(\mcsr/_0657_ ) );
OAI21_X1 \mcsr/_1534_ ( .A(\mcsr/_0657_ ), .B1(\mcsr/_0647_ ), .B2(\mcsr/_0556_ ), .ZN(\mcsr/_0849_ ) );
NAND4_X1 \mcsr/_1535_ ( .A1(\mcsr/_0654_ ), .A2(\mcsr/_0649_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0176_ ), .ZN(\mcsr/_0658_ ) );
OAI21_X1 \mcsr/_1536_ ( .A(\mcsr/_0658_ ), .B1(\mcsr/_0647_ ), .B2(\mcsr/_0563_ ), .ZN(\mcsr/_0850_ ) );
NAND4_X1 \mcsr/_1537_ ( .A1(\mcsr/_0654_ ), .A2(\mcsr/_0649_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0177_ ), .ZN(\mcsr/_0659_ ) );
OAI21_X1 \mcsr/_1538_ ( .A(\mcsr/_0659_ ), .B1(\mcsr/_0626_ ), .B2(\mcsr/_0570_ ), .ZN(\mcsr/_0851_ ) );
NAND4_X1 \mcsr/_1539_ ( .A1(\mcsr/_0654_ ), .A2(\mcsr/_0649_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0178_ ), .ZN(\mcsr/_0660_ ) );
OAI21_X1 \mcsr/_1540_ ( .A(\mcsr/_0660_ ), .B1(\mcsr/_0626_ ), .B2(\mcsr/_0577_ ), .ZN(\mcsr/_0852_ ) );
NAND4_X1 \mcsr/_1541_ ( .A1(\mcsr/_0654_ ), .A2(\mcsr/_0616_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0179_ ), .ZN(\mcsr/_0661_ ) );
OAI21_X1 \mcsr/_1542_ ( .A(\mcsr/_0661_ ), .B1(\mcsr/_0626_ ), .B2(\mcsr/_0584_ ), .ZN(\mcsr/_0853_ ) );
NAND4_X1 \mcsr/_1543_ ( .A1(\mcsr/_0654_ ), .A2(\mcsr/_0616_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0180_ ), .ZN(\mcsr/_0662_ ) );
OAI21_X1 \mcsr/_1544_ ( .A(\mcsr/_0662_ ), .B1(\mcsr/_0626_ ), .B2(\mcsr/_0591_ ), .ZN(\mcsr/_0854_ ) );
NAND4_X1 \mcsr/_1545_ ( .A1(\mcsr/_0654_ ), .A2(\mcsr/_0616_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0181_ ), .ZN(\mcsr/_0663_ ) );
OAI21_X1 \mcsr/_1546_ ( .A(\mcsr/_0663_ ), .B1(\mcsr/_0626_ ), .B2(\mcsr/_0598_ ), .ZN(\mcsr/_0855_ ) );
NAND4_X1 \mcsr/_1547_ ( .A1(\mcsr/_0654_ ), .A2(\mcsr/_0616_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0183_ ), .ZN(\mcsr/_0664_ ) );
OAI21_X1 \mcsr/_1548_ ( .A(\mcsr/_0664_ ), .B1(\mcsr/_0626_ ), .B2(\mcsr/_0605_ ), .ZN(\mcsr/_0857_ ) );
NAND4_X1 \mcsr/_1549_ ( .A1(\mcsr/_0619_ ), .A2(\mcsr/_0616_ ), .A3(\mcsr/_0269_ ), .A4(\mcsr/_0184_ ), .ZN(\mcsr/_0665_ ) );
OAI21_X1 \mcsr/_1550_ ( .A(\mcsr/_0665_ ), .B1(\mcsr/_0626_ ), .B2(\mcsr/_0612_ ), .ZN(\mcsr/_0858_ ) );
AND3_X2 \mcsr/_1551_ ( .A1(\mcsr/_0619_ ), .A2(\mcsr/_0898_ ), .A3(\mcsr/_0271_ ), .ZN(\mcsr/_0666_ ) );
NOR2_X1 \mcsr/_1552_ ( .A1(\mcsr/_0616_ ), .A2(\mcsr/_0269_ ), .ZN(\mcsr/_0667_ ) );
AND2_X1 \mcsr/_1553_ ( .A1(\mcsr/_0666_ ), .A2(\mcsr/_0667_ ), .ZN(\mcsr/_0668_ ) );
BUF_X4 \mcsr/_1554_ ( .A(\mcsr/_0668_ ), .Z(\mcsr/_0669_ ) );
AND2_X4 \mcsr/_1555_ ( .A1(\mcsr/_0369_ ), .A2(\mcsr/_0669_ ), .ZN(\mcsr/_0670_ ) );
BUF_X4 \mcsr/_1556_ ( .A(\mcsr/_0670_ ), .Z(\mcsr/_0671_ ) );
MUX2_X1 \mcsr/_1557_ ( .A(\mcsr/_0160_ ), .B(\mcsr/_0866_ ), .S(\mcsr/_0671_ ), .Z(\mcsr/_0000_ ) );
MUX2_X1 \mcsr/_1558_ ( .A(\mcsr/_0171_ ), .B(\mcsr/_0877_ ), .S(\mcsr/_0671_ ), .Z(\mcsr/_0001_ ) );
MUX2_X1 \mcsr/_1559_ ( .A(\mcsr/_0182_ ), .B(\mcsr/_0888_ ), .S(\mcsr/_0671_ ), .Z(\mcsr/_0002_ ) );
MUX2_X1 \mcsr/_1560_ ( .A(\mcsr/_0185_ ), .B(\mcsr/_0891_ ), .S(\mcsr/_0671_ ), .Z(\mcsr/_0003_ ) );
MUX2_X1 \mcsr/_1561_ ( .A(\mcsr/_0186_ ), .B(\mcsr/_0892_ ), .S(\mcsr/_0671_ ), .Z(\mcsr/_0004_ ) );
MUX2_X1 \mcsr/_1562_ ( .A(\mcsr/_0187_ ), .B(\mcsr/_0893_ ), .S(\mcsr/_0671_ ), .Z(\mcsr/_0005_ ) );
MUX2_X1 \mcsr/_1563_ ( .A(\mcsr/_0188_ ), .B(\mcsr/_0894_ ), .S(\mcsr/_0671_ ), .Z(\mcsr/_0006_ ) );
MUX2_X1 \mcsr/_1564_ ( .A(\mcsr/_0189_ ), .B(\mcsr/_0895_ ), .S(\mcsr/_0671_ ), .Z(\mcsr/_0007_ ) );
MUX2_X1 \mcsr/_1565_ ( .A(\mcsr/_0190_ ), .B(\mcsr/_0896_ ), .S(\mcsr/_0671_ ), .Z(\mcsr/_0008_ ) );
BUF_X4 \mcsr/_1566_ ( .A(\mcsr/_0670_ ), .Z(\mcsr/_0672_ ) );
MUX2_X1 \mcsr/_1567_ ( .A(\mcsr/_0191_ ), .B(\mcsr/_0897_ ), .S(\mcsr/_0672_ ), .Z(\mcsr/_0009_ ) );
MUX2_X1 \mcsr/_1568_ ( .A(\mcsr/_0161_ ), .B(\mcsr/_0867_ ), .S(\mcsr/_0672_ ), .Z(\mcsr/_0010_ ) );
INV_X1 \mcsr/_1569_ ( .A(\mcsr/_0669_ ), .ZN(\mcsr/_0673_ ) );
NOR3_X1 \mcsr/_1570_ ( .A1(\mcsr/_0371_ ), .A2(\mcsr/_0868_ ), .A3(\mcsr/_0673_ ), .ZN(\mcsr/_0674_ ) );
INV_X1 \mcsr/_1571_ ( .A(\mcsr/_0671_ ), .ZN(\mcsr/_0675_ ) );
AOI21_X1 \mcsr/_1572_ ( .A(\mcsr/_0674_ ), .B1(\mcsr/_0465_ ), .B2(\mcsr/_0675_ ), .ZN(\mcsr/_0011_ ) );
NOR3_X1 \mcsr/_1573_ ( .A1(\mcsr/_0371_ ), .A2(\mcsr/_0869_ ), .A3(\mcsr/_0673_ ), .ZN(\mcsr/_0676_ ) );
AOI21_X1 \mcsr/_1574_ ( .A(\mcsr/_0676_ ), .B1(\mcsr/_0470_ ), .B2(\mcsr/_0675_ ), .ZN(\mcsr/_0012_ ) );
MUX2_X1 \mcsr/_1575_ ( .A(\mcsr/_0164_ ), .B(\mcsr/_0870_ ), .S(\mcsr/_0672_ ), .Z(\mcsr/_0013_ ) );
MUX2_X1 \mcsr/_1576_ ( .A(\mcsr/_0165_ ), .B(\mcsr/_0871_ ), .S(\mcsr/_0672_ ), .Z(\mcsr/_0014_ ) );
MUX2_X1 \mcsr/_1577_ ( .A(\mcsr/_0166_ ), .B(\mcsr/_0872_ ), .S(\mcsr/_0672_ ), .Z(\mcsr/_0015_ ) );
MUX2_X1 \mcsr/_1578_ ( .A(\mcsr/_0167_ ), .B(\mcsr/_0873_ ), .S(\mcsr/_0672_ ), .Z(\mcsr/_0016_ ) );
MUX2_X1 \mcsr/_1579_ ( .A(\mcsr/_0168_ ), .B(\mcsr/_0874_ ), .S(\mcsr/_0672_ ), .Z(\mcsr/_0017_ ) );
MUX2_X1 \mcsr/_1580_ ( .A(\mcsr/_0169_ ), .B(\mcsr/_0875_ ), .S(\mcsr/_0672_ ), .Z(\mcsr/_0018_ ) );
MUX2_X1 \mcsr/_1581_ ( .A(\mcsr/_0170_ ), .B(\mcsr/_0876_ ), .S(\mcsr/_0672_ ), .Z(\mcsr/_0019_ ) );
MUX2_X1 \mcsr/_1582_ ( .A(\mcsr/_0172_ ), .B(\mcsr/_0878_ ), .S(\mcsr/_0672_ ), .Z(\mcsr/_0020_ ) );
BUF_X4 \mcsr/_1583_ ( .A(\mcsr/_0670_ ), .Z(\mcsr/_0677_ ) );
MUX2_X1 \mcsr/_1584_ ( .A(\mcsr/_0173_ ), .B(\mcsr/_0879_ ), .S(\mcsr/_0677_ ), .Z(\mcsr/_0021_ ) );
MUX2_X1 \mcsr/_1585_ ( .A(\mcsr/_0174_ ), .B(\mcsr/_0880_ ), .S(\mcsr/_0677_ ), .Z(\mcsr/_0022_ ) );
MUX2_X1 \mcsr/_1586_ ( .A(\mcsr/_0175_ ), .B(\mcsr/_0881_ ), .S(\mcsr/_0677_ ), .Z(\mcsr/_0023_ ) );
MUX2_X1 \mcsr/_1587_ ( .A(\mcsr/_0176_ ), .B(\mcsr/_0882_ ), .S(\mcsr/_0677_ ), .Z(\mcsr/_0024_ ) );
MUX2_X1 \mcsr/_1588_ ( .A(\mcsr/_0177_ ), .B(\mcsr/_0883_ ), .S(\mcsr/_0677_ ), .Z(\mcsr/_0025_ ) );
MUX2_X1 \mcsr/_1589_ ( .A(\mcsr/_0178_ ), .B(\mcsr/_0884_ ), .S(\mcsr/_0677_ ), .Z(\mcsr/_0026_ ) );
MUX2_X1 \mcsr/_1590_ ( .A(\mcsr/_0179_ ), .B(\mcsr/_0885_ ), .S(\mcsr/_0677_ ), .Z(\mcsr/_0027_ ) );
MUX2_X1 \mcsr/_1591_ ( .A(\mcsr/_0180_ ), .B(\mcsr/_0886_ ), .S(\mcsr/_0677_ ), .Z(\mcsr/_0028_ ) );
MUX2_X1 \mcsr/_1592_ ( .A(\mcsr/_0181_ ), .B(\mcsr/_0887_ ), .S(\mcsr/_0677_ ), .Z(\mcsr/_0029_ ) );
MUX2_X1 \mcsr/_1593_ ( .A(\mcsr/_0183_ ), .B(\mcsr/_0889_ ), .S(\mcsr/_0677_ ), .Z(\mcsr/_0030_ ) );
MUX2_X1 \mcsr/_1594_ ( .A(\mcsr/_0184_ ), .B(\mcsr/_0890_ ), .S(\mcsr/_0670_ ), .Z(\mcsr/_0031_ ) );
AND2_X4 \mcsr/_1595_ ( .A1(\mcsr/_0666_ ), .A2(\mcsr/_0640_ ), .ZN(\mcsr/_0678_ ) );
BUF_X4 \mcsr/_1596_ ( .A(\mcsr/_0678_ ), .Z(\mcsr/_0679_ ) );
MUX2_X1 \mcsr/_1597_ ( .A(\mcsr/_0866_ ), .B(\mcsr/_0770_ ), .S(\mcsr/_0679_ ), .Z(\mcsr/_0680_ ) );
NAND4_X1 \mcsr/_1598_ ( .A1(\mcsr/_0668_ ), .A2(\mcsr/_0355_ ), .A3(\mcsr/_0336_ ), .A4(\mcsr/_0458_ ), .ZN(\mcsr/_0681_ ) );
INV_X2 \mcsr/_1599_ ( .A(\mcsr/_0678_ ), .ZN(\mcsr/_0682_ ) );
AND2_X4 \mcsr/_1600_ ( .A1(\mcsr/_0681_ ), .A2(\mcsr/_0682_ ), .ZN(\mcsr/_0683_ ) );
BUF_X4 \mcsr/_1601_ ( .A(\mcsr/_0683_ ), .Z(\mcsr/_0684_ ) );
MUX2_X1 \mcsr/_1602_ ( .A(\mcsr/_0680_ ), .B(\mcsr/_0192_ ), .S(\mcsr/_0684_ ), .Z(\mcsr/_0032_ ) );
MUX2_X1 \mcsr/_1603_ ( .A(\mcsr/_0877_ ), .B(\mcsr/_0781_ ), .S(\mcsr/_0679_ ), .Z(\mcsr/_0685_ ) );
MUX2_X1 \mcsr/_1604_ ( .A(\mcsr/_0685_ ), .B(\mcsr/_0203_ ), .S(\mcsr/_0684_ ), .Z(\mcsr/_0033_ ) );
BUF_X4 \mcsr/_1605_ ( .A(\mcsr/_0682_ ), .Z(\mcsr/_0686_ ) );
NAND2_X1 \mcsr/_1606_ ( .A1(\mcsr/_0345_ ), .A2(\mcsr/_0669_ ), .ZN(\mcsr/_0687_ ) );
BUF_X4 \mcsr/_1607_ ( .A(\mcsr/_0687_ ), .Z(\mcsr/_0688_ ) );
OAI21_X1 \mcsr/_1608_ ( .A(\mcsr/_0686_ ), .B1(\mcsr/_0688_ ), .B2(\mcsr/_0888_ ), .ZN(\mcsr/_0689_ ) );
BUF_X4 \mcsr/_1609_ ( .A(\mcsr/_0666_ ), .Z(\mcsr/_0690_ ) );
NAND3_X1 \mcsr/_1610_ ( .A1(\mcsr/_0690_ ), .A2(\mcsr/_0792_ ), .A3(\mcsr/_0641_ ), .ZN(\mcsr/_0691_ ) );
BUF_X4 \mcsr/_1611_ ( .A(\mcsr/_0683_ ), .Z(\mcsr/_0692_ ) );
AOI22_X1 \mcsr/_1612_ ( .A1(\mcsr/_0689_ ), .A2(\mcsr/_0691_ ), .B1(\mcsr/_0692_ ), .B2(\mcsr/_0389_ ), .ZN(\mcsr/_0034_ ) );
MUX2_X1 \mcsr/_1613_ ( .A(\mcsr/_0891_ ), .B(\mcsr/_0795_ ), .S(\mcsr/_0679_ ), .Z(\mcsr/_0693_ ) );
MUX2_X1 \mcsr/_1614_ ( .A(\mcsr/_0693_ ), .B(\mcsr/_0217_ ), .S(\mcsr/_0684_ ), .Z(\mcsr/_0035_ ) );
MUX2_X1 \mcsr/_1615_ ( .A(\mcsr/_0892_ ), .B(\mcsr/_0796_ ), .S(\mcsr/_0679_ ), .Z(\mcsr/_0694_ ) );
MUX2_X1 \mcsr/_1616_ ( .A(\mcsr/_0694_ ), .B(\mcsr/_0218_ ), .S(\mcsr/_0684_ ), .Z(\mcsr/_0036_ ) );
MUX2_X1 \mcsr/_1617_ ( .A(\mcsr/_0893_ ), .B(\mcsr/_0797_ ), .S(\mcsr/_0679_ ), .Z(\mcsr/_0695_ ) );
MUX2_X1 \mcsr/_1618_ ( .A(\mcsr/_0695_ ), .B(\mcsr/_0219_ ), .S(\mcsr/_0684_ ), .Z(\mcsr/_0037_ ) );
MUX2_X1 \mcsr/_1619_ ( .A(\mcsr/_0894_ ), .B(\mcsr/_0798_ ), .S(\mcsr/_0679_ ), .Z(\mcsr/_0696_ ) );
MUX2_X1 \mcsr/_1620_ ( .A(\mcsr/_0696_ ), .B(\mcsr/_0220_ ), .S(\mcsr/_0684_ ), .Z(\mcsr/_0038_ ) );
MUX2_X1 \mcsr/_1621_ ( .A(\mcsr/_0895_ ), .B(\mcsr/_0799_ ), .S(\mcsr/_0679_ ), .Z(\mcsr/_0697_ ) );
MUX2_X1 \mcsr/_1622_ ( .A(\mcsr/_0697_ ), .B(\mcsr/_0221_ ), .S(\mcsr/_0684_ ), .Z(\mcsr/_0039_ ) );
OAI21_X1 \mcsr/_1623_ ( .A(\mcsr/_0686_ ), .B1(\mcsr/_0688_ ), .B2(\mcsr/_0896_ ), .ZN(\mcsr/_0698_ ) );
NAND3_X1 \mcsr/_1624_ ( .A1(\mcsr/_0690_ ), .A2(\mcsr/_0800_ ), .A3(\mcsr/_0641_ ), .ZN(\mcsr/_0699_ ) );
AOI22_X1 \mcsr/_1625_ ( .A1(\mcsr/_0698_ ), .A2(\mcsr/_0699_ ), .B1(\mcsr/_0692_ ), .B2(\mcsr/_0437_ ), .ZN(\mcsr/_0040_ ) );
OAI21_X1 \mcsr/_1626_ ( .A(\mcsr/_0686_ ), .B1(\mcsr/_0688_ ), .B2(\mcsr/_0897_ ), .ZN(\mcsr/_0700_ ) );
NAND3_X1 \mcsr/_1627_ ( .A1(\mcsr/_0690_ ), .A2(\mcsr/_0801_ ), .A3(\mcsr/_0641_ ), .ZN(\mcsr/_0701_ ) );
AOI22_X1 \mcsr/_1628_ ( .A1(\mcsr/_0700_ ), .A2(\mcsr/_0701_ ), .B1(\mcsr/_0692_ ), .B2(\mcsr/_0446_ ), .ZN(\mcsr/_0041_ ) );
OAI21_X1 \mcsr/_1629_ ( .A(\mcsr/_0686_ ), .B1(\mcsr/_0688_ ), .B2(\mcsr/_0867_ ), .ZN(\mcsr/_0702_ ) );
NAND3_X1 \mcsr/_1630_ ( .A1(\mcsr/_0690_ ), .A2(\mcsr/_0771_ ), .A3(\mcsr/_0641_ ), .ZN(\mcsr/_0703_ ) );
AOI22_X1 \mcsr/_1631_ ( .A1(\mcsr/_0702_ ), .A2(\mcsr/_0703_ ), .B1(\mcsr/_0692_ ), .B2(\mcsr/_0453_ ), .ZN(\mcsr/_0042_ ) );
MUX2_X1 \mcsr/_1632_ ( .A(\mcsr/_0868_ ), .B(\mcsr/_0772_ ), .S(\mcsr/_0679_ ), .Z(\mcsr/_0704_ ) );
MUX2_X1 \mcsr/_1633_ ( .A(\mcsr/_0704_ ), .B(\mcsr/_0194_ ), .S(\mcsr/_0683_ ), .Z(\mcsr/_0043_ ) );
MUX2_X1 \mcsr/_1634_ ( .A(\mcsr/_0869_ ), .B(\mcsr/_0773_ ), .S(\mcsr/_0678_ ), .Z(\mcsr/_0705_ ) );
MUX2_X1 \mcsr/_1635_ ( .A(\mcsr/_0705_ ), .B(\mcsr/_0195_ ), .S(\mcsr/_0683_ ), .Z(\mcsr/_0044_ ) );
OAI21_X1 \mcsr/_1636_ ( .A(\mcsr/_0686_ ), .B1(\mcsr/_0688_ ), .B2(\mcsr/_0870_ ), .ZN(\mcsr/_0706_ ) );
NAND3_X1 \mcsr/_1637_ ( .A1(\mcsr/_0690_ ), .A2(\mcsr/_0774_ ), .A3(\mcsr/_0641_ ), .ZN(\mcsr/_0707_ ) );
AOI22_X1 \mcsr/_1638_ ( .A1(\mcsr/_0706_ ), .A2(\mcsr/_0707_ ), .B1(\mcsr/_0692_ ), .B2(\mcsr/_0478_ ), .ZN(\mcsr/_0045_ ) );
OAI21_X1 \mcsr/_1639_ ( .A(\mcsr/_0686_ ), .B1(\mcsr/_0688_ ), .B2(\mcsr/_0871_ ), .ZN(\mcsr/_0708_ ) );
NAND3_X1 \mcsr/_1640_ ( .A1(\mcsr/_0690_ ), .A2(\mcsr/_0775_ ), .A3(\mcsr/_0641_ ), .ZN(\mcsr/_0709_ ) );
AOI22_X1 \mcsr/_1641_ ( .A1(\mcsr/_0708_ ), .A2(\mcsr/_0709_ ), .B1(\mcsr/_0692_ ), .B2(\mcsr/_0485_ ), .ZN(\mcsr/_0046_ ) );
OAI21_X1 \mcsr/_1642_ ( .A(\mcsr/_0686_ ), .B1(\mcsr/_0688_ ), .B2(\mcsr/_0872_ ), .ZN(\mcsr/_0710_ ) );
NAND3_X1 \mcsr/_1643_ ( .A1(\mcsr/_0690_ ), .A2(\mcsr/_0776_ ), .A3(\mcsr/_0641_ ), .ZN(\mcsr/_0711_ ) );
AOI22_X1 \mcsr/_1644_ ( .A1(\mcsr/_0710_ ), .A2(\mcsr/_0711_ ), .B1(\mcsr/_0692_ ), .B2(\mcsr/_0493_ ), .ZN(\mcsr/_0047_ ) );
BUF_X4 \mcsr/_1645_ ( .A(\mcsr/_0682_ ), .Z(\mcsr/_0712_ ) );
OAI21_X1 \mcsr/_1646_ ( .A(\mcsr/_0712_ ), .B1(\mcsr/_0688_ ), .B2(\mcsr/_0873_ ), .ZN(\mcsr/_0713_ ) );
NAND3_X1 \mcsr/_1647_ ( .A1(\mcsr/_0690_ ), .A2(\mcsr/_0777_ ), .A3(\mcsr/_0641_ ), .ZN(\mcsr/_0714_ ) );
AOI22_X1 \mcsr/_1648_ ( .A1(\mcsr/_0713_ ), .A2(\mcsr/_0714_ ), .B1(\mcsr/_0692_ ), .B2(\mcsr/_0504_ ), .ZN(\mcsr/_0048_ ) );
OAI21_X1 \mcsr/_1649_ ( .A(\mcsr/_0712_ ), .B1(\mcsr/_0688_ ), .B2(\mcsr/_0874_ ), .ZN(\mcsr/_0715_ ) );
NAND3_X1 \mcsr/_1650_ ( .A1(\mcsr/_0690_ ), .A2(\mcsr/_0778_ ), .A3(\mcsr/_0641_ ), .ZN(\mcsr/_0716_ ) );
AOI22_X1 \mcsr/_1651_ ( .A1(\mcsr/_0715_ ), .A2(\mcsr/_0716_ ), .B1(\mcsr/_0692_ ), .B2(\mcsr/_0511_ ), .ZN(\mcsr/_0049_ ) );
OAI21_X1 \mcsr/_1652_ ( .A(\mcsr/_0712_ ), .B1(\mcsr/_0688_ ), .B2(\mcsr/_0875_ ), .ZN(\mcsr/_0717_ ) );
BUF_X4 \mcsr/_1653_ ( .A(\mcsr/_0640_ ), .Z(\mcsr/_0718_ ) );
NAND3_X1 \mcsr/_1654_ ( .A1(\mcsr/_0690_ ), .A2(\mcsr/_0779_ ), .A3(\mcsr/_0718_ ), .ZN(\mcsr/_0719_ ) );
AOI22_X1 \mcsr/_1655_ ( .A1(\mcsr/_0717_ ), .A2(\mcsr/_0719_ ), .B1(\mcsr/_0692_ ), .B2(\mcsr/_0519_ ), .ZN(\mcsr/_0050_ ) );
BUF_X4 \mcsr/_1656_ ( .A(\mcsr/_0687_ ), .Z(\mcsr/_0720_ ) );
OAI21_X1 \mcsr/_1657_ ( .A(\mcsr/_0712_ ), .B1(\mcsr/_0720_ ), .B2(\mcsr/_0876_ ), .ZN(\mcsr/_0721_ ) );
BUF_X4 \mcsr/_1658_ ( .A(\mcsr/_0666_ ), .Z(\mcsr/_0722_ ) );
NAND3_X1 \mcsr/_1659_ ( .A1(\mcsr/_0722_ ), .A2(\mcsr/_0780_ ), .A3(\mcsr/_0718_ ), .ZN(\mcsr/_0723_ ) );
BUF_X4 \mcsr/_1660_ ( .A(\mcsr/_0683_ ), .Z(\mcsr/_0724_ ) );
AOI22_X1 \mcsr/_1661_ ( .A1(\mcsr/_0721_ ), .A2(\mcsr/_0723_ ), .B1(\mcsr/_0724_ ), .B2(\mcsr/_0526_ ), .ZN(\mcsr/_0051_ ) );
OAI21_X1 \mcsr/_1662_ ( .A(\mcsr/_0712_ ), .B1(\mcsr/_0720_ ), .B2(\mcsr/_0878_ ), .ZN(\mcsr/_0725_ ) );
NAND3_X1 \mcsr/_1663_ ( .A1(\mcsr/_0722_ ), .A2(\mcsr/_0782_ ), .A3(\mcsr/_0718_ ), .ZN(\mcsr/_0726_ ) );
AOI22_X1 \mcsr/_1664_ ( .A1(\mcsr/_0725_ ), .A2(\mcsr/_0726_ ), .B1(\mcsr/_0724_ ), .B2(\mcsr/_0533_ ), .ZN(\mcsr/_0052_ ) );
OAI21_X1 \mcsr/_1665_ ( .A(\mcsr/_0712_ ), .B1(\mcsr/_0720_ ), .B2(\mcsr/_0879_ ), .ZN(\mcsr/_0727_ ) );
NAND3_X1 \mcsr/_1666_ ( .A1(\mcsr/_0722_ ), .A2(\mcsr/_0783_ ), .A3(\mcsr/_0718_ ), .ZN(\mcsr/_0728_ ) );
AOI22_X1 \mcsr/_1667_ ( .A1(\mcsr/_0727_ ), .A2(\mcsr/_0728_ ), .B1(\mcsr/_0724_ ), .B2(\mcsr/_0542_ ), .ZN(\mcsr/_0053_ ) );
OAI21_X1 \mcsr/_1668_ ( .A(\mcsr/_0712_ ), .B1(\mcsr/_0720_ ), .B2(\mcsr/_0880_ ), .ZN(\mcsr/_0729_ ) );
NAND3_X1 \mcsr/_1669_ ( .A1(\mcsr/_0722_ ), .A2(\mcsr/_0784_ ), .A3(\mcsr/_0718_ ), .ZN(\mcsr/_0730_ ) );
AOI22_X1 \mcsr/_1670_ ( .A1(\mcsr/_0729_ ), .A2(\mcsr/_0730_ ), .B1(\mcsr/_0724_ ), .B2(\mcsr/_0549_ ), .ZN(\mcsr/_0054_ ) );
OAI21_X1 \mcsr/_1671_ ( .A(\mcsr/_0712_ ), .B1(\mcsr/_0720_ ), .B2(\mcsr/_0881_ ), .ZN(\mcsr/_0731_ ) );
NAND3_X1 \mcsr/_1672_ ( .A1(\mcsr/_0722_ ), .A2(\mcsr/_0785_ ), .A3(\mcsr/_0718_ ), .ZN(\mcsr/_0732_ ) );
AOI22_X1 \mcsr/_1673_ ( .A1(\mcsr/_0731_ ), .A2(\mcsr/_0732_ ), .B1(\mcsr/_0724_ ), .B2(\mcsr/_0556_ ), .ZN(\mcsr/_0055_ ) );
OAI21_X1 \mcsr/_1674_ ( .A(\mcsr/_0712_ ), .B1(\mcsr/_0720_ ), .B2(\mcsr/_0882_ ), .ZN(\mcsr/_0733_ ) );
NAND3_X1 \mcsr/_1675_ ( .A1(\mcsr/_0722_ ), .A2(\mcsr/_0786_ ), .A3(\mcsr/_0718_ ), .ZN(\mcsr/_0734_ ) );
AOI22_X1 \mcsr/_1676_ ( .A1(\mcsr/_0733_ ), .A2(\mcsr/_0734_ ), .B1(\mcsr/_0724_ ), .B2(\mcsr/_0563_ ), .ZN(\mcsr/_0056_ ) );
OAI21_X1 \mcsr/_1677_ ( .A(\mcsr/_0712_ ), .B1(\mcsr/_0720_ ), .B2(\mcsr/_0883_ ), .ZN(\mcsr/_0735_ ) );
NAND3_X1 \mcsr/_1678_ ( .A1(\mcsr/_0722_ ), .A2(\mcsr/_0787_ ), .A3(\mcsr/_0718_ ), .ZN(\mcsr/_0736_ ) );
AOI22_X1 \mcsr/_1679_ ( .A1(\mcsr/_0735_ ), .A2(\mcsr/_0736_ ), .B1(\mcsr/_0724_ ), .B2(\mcsr/_0570_ ), .ZN(\mcsr/_0057_ ) );
OAI21_X1 \mcsr/_1680_ ( .A(\mcsr/_0682_ ), .B1(\mcsr/_0720_ ), .B2(\mcsr/_0884_ ), .ZN(\mcsr/_0737_ ) );
NAND3_X1 \mcsr/_1681_ ( .A1(\mcsr/_0722_ ), .A2(\mcsr/_0788_ ), .A3(\mcsr/_0718_ ), .ZN(\mcsr/_0738_ ) );
AOI22_X1 \mcsr/_1682_ ( .A1(\mcsr/_0737_ ), .A2(\mcsr/_0738_ ), .B1(\mcsr/_0724_ ), .B2(\mcsr/_0577_ ), .ZN(\mcsr/_0058_ ) );
OAI21_X1 \mcsr/_1683_ ( .A(\mcsr/_0682_ ), .B1(\mcsr/_0720_ ), .B2(\mcsr/_0885_ ), .ZN(\mcsr/_0739_ ) );
NAND3_X1 \mcsr/_1684_ ( .A1(\mcsr/_0722_ ), .A2(\mcsr/_0789_ ), .A3(\mcsr/_0718_ ), .ZN(\mcsr/_0740_ ) );
AOI22_X1 \mcsr/_1685_ ( .A1(\mcsr/_0739_ ), .A2(\mcsr/_0740_ ), .B1(\mcsr/_0724_ ), .B2(\mcsr/_0584_ ), .ZN(\mcsr/_0059_ ) );
OAI21_X1 \mcsr/_1686_ ( .A(\mcsr/_0682_ ), .B1(\mcsr/_0720_ ), .B2(\mcsr/_0886_ ), .ZN(\mcsr/_0741_ ) );
NAND3_X1 \mcsr/_1687_ ( .A1(\mcsr/_0722_ ), .A2(\mcsr/_0790_ ), .A3(\mcsr/_0640_ ), .ZN(\mcsr/_0742_ ) );
AOI22_X1 \mcsr/_1688_ ( .A1(\mcsr/_0741_ ), .A2(\mcsr/_0742_ ), .B1(\mcsr/_0724_ ), .B2(\mcsr/_0591_ ), .ZN(\mcsr/_0060_ ) );
OAI21_X1 \mcsr/_1689_ ( .A(\mcsr/_0682_ ), .B1(\mcsr/_0687_ ), .B2(\mcsr/_0887_ ), .ZN(\mcsr/_0743_ ) );
NAND3_X1 \mcsr/_1690_ ( .A1(\mcsr/_0666_ ), .A2(\mcsr/_0791_ ), .A3(\mcsr/_0640_ ), .ZN(\mcsr/_0744_ ) );
AOI22_X1 \mcsr/_1691_ ( .A1(\mcsr/_0743_ ), .A2(\mcsr/_0744_ ), .B1(\mcsr/_0684_ ), .B2(\mcsr/_0598_ ), .ZN(\mcsr/_0061_ ) );
OAI21_X1 \mcsr/_1692_ ( .A(\mcsr/_0682_ ), .B1(\mcsr/_0687_ ), .B2(\mcsr/_0889_ ), .ZN(\mcsr/_0745_ ) );
NAND3_X1 \mcsr/_1693_ ( .A1(\mcsr/_0666_ ), .A2(\mcsr/_0793_ ), .A3(\mcsr/_0640_ ), .ZN(\mcsr/_0746_ ) );
AOI22_X1 \mcsr/_1694_ ( .A1(\mcsr/_0745_ ), .A2(\mcsr/_0746_ ), .B1(\mcsr/_0684_ ), .B2(\mcsr/_0605_ ), .ZN(\mcsr/_0062_ ) );
OAI21_X1 \mcsr/_1695_ ( .A(\mcsr/_0682_ ), .B1(\mcsr/_0687_ ), .B2(\mcsr/_0890_ ), .ZN(\mcsr/_0747_ ) );
NAND3_X1 \mcsr/_1696_ ( .A1(\mcsr/_0666_ ), .A2(\mcsr/_0794_ ), .A3(\mcsr/_0640_ ), .ZN(\mcsr/_0748_ ) );
AOI22_X1 \mcsr/_1697_ ( .A1(\mcsr/_0747_ ), .A2(\mcsr/_0748_ ), .B1(\mcsr/_0684_ ), .B2(\mcsr/_0612_ ), .ZN(\mcsr/_0063_ ) );
NOR3_X1 \mcsr/_1698_ ( .A1(\mcsr/_0342_ ), .A2(\mcsr/_0345_ ), .A3(\mcsr/_0369_ ), .ZN(\mcsr/_0749_ ) );
NAND2_X2 \mcsr/_1699_ ( .A1(\mcsr/_0749_ ), .A2(\mcsr/_0668_ ), .ZN(\mcsr/_0750_ ) );
BUF_X4 \mcsr/_1700_ ( .A(\mcsr/_0750_ ), .Z(\mcsr/_0751_ ) );
MUX2_X1 \mcsr/_1701_ ( .A(\mcsr/_0866_ ), .B(\mcsr/_0128_ ), .S(\mcsr/_0751_ ), .Z(\mcsr/_0096_ ) );
MUX2_X1 \mcsr/_1702_ ( .A(\mcsr/_0877_ ), .B(\mcsr/_0139_ ), .S(\mcsr/_0751_ ), .Z(\mcsr/_0097_ ) );
MUX2_X1 \mcsr/_1703_ ( .A(\mcsr/_0888_ ), .B(\mcsr/_0150_ ), .S(\mcsr/_0751_ ), .Z(\mcsr/_0098_ ) );
MUX2_X1 \mcsr/_1704_ ( .A(\mcsr/_0891_ ), .B(\mcsr/_0153_ ), .S(\mcsr/_0751_ ), .Z(\mcsr/_0099_ ) );
MUX2_X1 \mcsr/_1705_ ( .A(\mcsr/_0892_ ), .B(\mcsr/_0154_ ), .S(\mcsr/_0751_ ), .Z(\mcsr/_0100_ ) );
MUX2_X1 \mcsr/_1706_ ( .A(\mcsr/_0893_ ), .B(\mcsr/_0155_ ), .S(\mcsr/_0751_ ), .Z(\mcsr/_0101_ ) );
MUX2_X1 \mcsr/_1707_ ( .A(\mcsr/_0894_ ), .B(\mcsr/_0156_ ), .S(\mcsr/_0751_ ), .Z(\mcsr/_0102_ ) );
MUX2_X1 \mcsr/_1708_ ( .A(\mcsr/_0895_ ), .B(\mcsr/_0157_ ), .S(\mcsr/_0751_ ), .Z(\mcsr/_0103_ ) );
MUX2_X1 \mcsr/_1709_ ( .A(\mcsr/_0896_ ), .B(\mcsr/_0158_ ), .S(\mcsr/_0751_ ), .Z(\mcsr/_0104_ ) );
MUX2_X1 \mcsr/_1710_ ( .A(\mcsr/_0897_ ), .B(\mcsr/_0159_ ), .S(\mcsr/_0751_ ), .Z(\mcsr/_0105_ ) );
BUF_X4 \mcsr/_1711_ ( .A(\mcsr/_0750_ ), .Z(\mcsr/_0752_ ) );
MUX2_X1 \mcsr/_1712_ ( .A(\mcsr/_0867_ ), .B(\mcsr/_0129_ ), .S(\mcsr/_0752_ ), .Z(\mcsr/_0106_ ) );
MUX2_X1 \mcsr/_1713_ ( .A(\mcsr/_0868_ ), .B(\mcsr/_0130_ ), .S(\mcsr/_0752_ ), .Z(\mcsr/_0107_ ) );
MUX2_X1 \mcsr/_1714_ ( .A(\mcsr/_0869_ ), .B(\mcsr/_0131_ ), .S(\mcsr/_0752_ ), .Z(\mcsr/_0108_ ) );
MUX2_X1 \mcsr/_1715_ ( .A(\mcsr/_0870_ ), .B(\mcsr/_0132_ ), .S(\mcsr/_0752_ ), .Z(\mcsr/_0109_ ) );
MUX2_X1 \mcsr/_1716_ ( .A(\mcsr/_0871_ ), .B(\mcsr/_0133_ ), .S(\mcsr/_0752_ ), .Z(\mcsr/_0110_ ) );
MUX2_X1 \mcsr/_1717_ ( .A(\mcsr/_0872_ ), .B(\mcsr/_0134_ ), .S(\mcsr/_0752_ ), .Z(\mcsr/_0111_ ) );
MUX2_X1 \mcsr/_1718_ ( .A(\mcsr/_0873_ ), .B(\mcsr/_0135_ ), .S(\mcsr/_0752_ ), .Z(\mcsr/_0112_ ) );
MUX2_X1 \mcsr/_1719_ ( .A(\mcsr/_0874_ ), .B(\mcsr/_0136_ ), .S(\mcsr/_0752_ ), .Z(\mcsr/_0113_ ) );
MUX2_X1 \mcsr/_1720_ ( .A(\mcsr/_0875_ ), .B(\mcsr/_0137_ ), .S(\mcsr/_0752_ ), .Z(\mcsr/_0114_ ) );
MUX2_X1 \mcsr/_1721_ ( .A(\mcsr/_0876_ ), .B(\mcsr/_0138_ ), .S(\mcsr/_0752_ ), .Z(\mcsr/_0115_ ) );
BUF_X4 \mcsr/_1722_ ( .A(\mcsr/_0750_ ), .Z(\mcsr/_0753_ ) );
MUX2_X1 \mcsr/_1723_ ( .A(\mcsr/_0878_ ), .B(\mcsr/_0140_ ), .S(\mcsr/_0753_ ), .Z(\mcsr/_0116_ ) );
MUX2_X1 \mcsr/_1724_ ( .A(\mcsr/_0879_ ), .B(\mcsr/_0141_ ), .S(\mcsr/_0753_ ), .Z(\mcsr/_0117_ ) );
MUX2_X1 \mcsr/_1725_ ( .A(\mcsr/_0880_ ), .B(\mcsr/_0142_ ), .S(\mcsr/_0753_ ), .Z(\mcsr/_0118_ ) );
MUX2_X1 \mcsr/_1726_ ( .A(\mcsr/_0881_ ), .B(\mcsr/_0143_ ), .S(\mcsr/_0753_ ), .Z(\mcsr/_0119_ ) );
MUX2_X1 \mcsr/_1727_ ( .A(\mcsr/_0882_ ), .B(\mcsr/_0144_ ), .S(\mcsr/_0753_ ), .Z(\mcsr/_0120_ ) );
MUX2_X1 \mcsr/_1728_ ( .A(\mcsr/_0883_ ), .B(\mcsr/_0145_ ), .S(\mcsr/_0753_ ), .Z(\mcsr/_0121_ ) );
MUX2_X1 \mcsr/_1729_ ( .A(\mcsr/_0884_ ), .B(\mcsr/_0146_ ), .S(\mcsr/_0753_ ), .Z(\mcsr/_0122_ ) );
MUX2_X1 \mcsr/_1730_ ( .A(\mcsr/_0885_ ), .B(\mcsr/_0147_ ), .S(\mcsr/_0753_ ), .Z(\mcsr/_0123_ ) );
MUX2_X1 \mcsr/_1731_ ( .A(\mcsr/_0886_ ), .B(\mcsr/_0148_ ), .S(\mcsr/_0753_ ), .Z(\mcsr/_0124_ ) );
MUX2_X1 \mcsr/_1732_ ( .A(\mcsr/_0887_ ), .B(\mcsr/_0149_ ), .S(\mcsr/_0753_ ), .Z(\mcsr/_0125_ ) );
MUX2_X1 \mcsr/_1733_ ( .A(\mcsr/_0889_ ), .B(\mcsr/_0151_ ), .S(\mcsr/_0750_ ), .Z(\mcsr/_0126_ ) );
MUX2_X1 \mcsr/_1734_ ( .A(\mcsr/_0890_ ), .B(\mcsr/_0152_ ), .S(\mcsr/_0750_ ), .Z(\mcsr/_0127_ ) );
BUF_X4 \mcsr/_1735_ ( .A(\mcsr/_0339_ ), .Z(\mcsr/_0754_ ) );
BUF_X4 \mcsr/_1736_ ( .A(\mcsr/_0341_ ), .Z(\mcsr/_0755_ ) );
BUF_X4 \mcsr/_1737_ ( .A(\mcsr/_0669_ ), .Z(\mcsr/_0756_ ) );
NAND4_X1 \mcsr/_1738_ ( .A1(\mcsr/_0754_ ), .A2(\mcsr/_0866_ ), .A3(\mcsr/_0755_ ), .A4(\mcsr/_0756_ ), .ZN(\mcsr/_0757_ ) );
AND2_X2 \mcsr/_1739_ ( .A1(\mcsr/_0357_ ), .A2(\mcsr/_0669_ ), .ZN(\mcsr/_0758_ ) );
OAI211_X2 \mcsr/_1740_ ( .A(\mcsr/_0686_ ), .B(\mcsr/_0757_ ), .C1(\mcsr/_0758_ ), .C2(\mcsr/_0353_ ), .ZN(\mcsr/_0064_ ) );
NAND4_X1 \mcsr/_1741_ ( .A1(\mcsr/_0339_ ), .A2(\mcsr/_0877_ ), .A3(\mcsr/_0341_ ), .A4(\mcsr/_0669_ ), .ZN(\mcsr/_0759_ ) );
OAI211_X2 \mcsr/_1742_ ( .A(\mcsr/_0686_ ), .B(\mcsr/_0759_ ), .C1(\mcsr/_0758_ ), .C2(\mcsr/_0380_ ), .ZN(\mcsr/_0065_ ) );
BUF_X4 \mcsr/_1743_ ( .A(\mcsr/_0679_ ), .Z(\mcsr/_0760_ ) );
BUF_X4 \mcsr/_1744_ ( .A(\mcsr/_0760_ ), .Z(\mcsr/_0761_ ) );
NAND2_X1 \mcsr/_1745_ ( .A1(\mcsr/_0357_ ), .A2(\mcsr/_0669_ ), .ZN(\mcsr/_0762_ ) );
BUF_X4 \mcsr/_1746_ ( .A(\mcsr/_0762_ ), .Z(\mcsr/_0763_ ) );
BUF_X4 \mcsr/_1747_ ( .A(\mcsr/_0763_ ), .Z(\mcsr/_0764_ ) );
NAND2_X1 \mcsr/_1748_ ( .A1(\mcsr/_0764_ ), .A2(\mcsr/_0246_ ), .ZN(\mcsr/_0765_ ) );
BUF_X4 \mcsr/_1749_ ( .A(\mcsr/_0339_ ), .Z(\mcsr/_0766_ ) );
BUF_X4 \mcsr/_1750_ ( .A(\mcsr/_0341_ ), .Z(\mcsr/_0767_ ) );
BUF_X4 \mcsr/_1751_ ( .A(\mcsr/_0669_ ), .Z(\mcsr/_0768_ ) );
NAND4_X1 \mcsr/_1752_ ( .A1(\mcsr/_0766_ ), .A2(\mcsr/_0888_ ), .A3(\mcsr/_0767_ ), .A4(\mcsr/_0768_ ), .ZN(\mcsr/_0769_ ) );
AOI21_X1 \mcsr/_1753_ ( .A(\mcsr/_0761_ ), .B1(\mcsr/_0765_ ), .B2(\mcsr/_0769_ ), .ZN(\mcsr/_0066_ ) );
NAND4_X1 \mcsr/_1754_ ( .A1(\mcsr/_0339_ ), .A2(\mcsr/_0891_ ), .A3(\mcsr/_0341_ ), .A4(\mcsr/_0669_ ), .ZN(\mcsr/_0272_ ) );
OAI211_X2 \mcsr/_1755_ ( .A(\mcsr/_0686_ ), .B(\mcsr/_0272_ ), .C1(\mcsr/_0758_ ), .C2(\mcsr/_0399_ ), .ZN(\mcsr/_0067_ ) );
NAND2_X1 \mcsr/_1756_ ( .A1(\mcsr/_0764_ ), .A2(\mcsr/_0250_ ), .ZN(\mcsr/_0273_ ) );
NAND4_X1 \mcsr/_1757_ ( .A1(\mcsr/_0766_ ), .A2(\mcsr/_0892_ ), .A3(\mcsr/_0767_ ), .A4(\mcsr/_0768_ ), .ZN(\mcsr/_0274_ ) );
AOI21_X1 \mcsr/_1758_ ( .A(\mcsr/_0761_ ), .B1(\mcsr/_0273_ ), .B2(\mcsr/_0274_ ), .ZN(\mcsr/_0068_ ) );
NAND2_X1 \mcsr/_1759_ ( .A1(\mcsr/_0764_ ), .A2(\mcsr/_0251_ ), .ZN(\mcsr/_0275_ ) );
NAND4_X1 \mcsr/_1760_ ( .A1(\mcsr/_0766_ ), .A2(\mcsr/_0893_ ), .A3(\mcsr/_0767_ ), .A4(\mcsr/_0768_ ), .ZN(\mcsr/_0276_ ) );
AOI21_X1 \mcsr/_1761_ ( .A(\mcsr/_0761_ ), .B1(\mcsr/_0275_ ), .B2(\mcsr/_0276_ ), .ZN(\mcsr/_0069_ ) );
NAND2_X1 \mcsr/_1762_ ( .A1(\mcsr/_0764_ ), .A2(\mcsr/_0252_ ), .ZN(\mcsr/_0277_ ) );
NAND4_X1 \mcsr/_1763_ ( .A1(\mcsr/_0766_ ), .A2(\mcsr/_0894_ ), .A3(\mcsr/_0767_ ), .A4(\mcsr/_0768_ ), .ZN(\mcsr/_0278_ ) );
AOI21_X1 \mcsr/_1764_ ( .A(\mcsr/_0761_ ), .B1(\mcsr/_0277_ ), .B2(\mcsr/_0278_ ), .ZN(\mcsr/_0070_ ) );
NAND2_X1 \mcsr/_1765_ ( .A1(\mcsr/_0764_ ), .A2(\mcsr/_0253_ ), .ZN(\mcsr/_0279_ ) );
NAND4_X1 \mcsr/_1766_ ( .A1(\mcsr/_0766_ ), .A2(\mcsr/_0895_ ), .A3(\mcsr/_0767_ ), .A4(\mcsr/_0768_ ), .ZN(\mcsr/_0280_ ) );
AOI21_X1 \mcsr/_1767_ ( .A(\mcsr/_0761_ ), .B1(\mcsr/_0279_ ), .B2(\mcsr/_0280_ ), .ZN(\mcsr/_0071_ ) );
NAND2_X1 \mcsr/_1768_ ( .A1(\mcsr/_0764_ ), .A2(\mcsr/_0254_ ), .ZN(\mcsr/_0281_ ) );
NAND4_X1 \mcsr/_1769_ ( .A1(\mcsr/_0766_ ), .A2(\mcsr/_0896_ ), .A3(\mcsr/_0767_ ), .A4(\mcsr/_0768_ ), .ZN(\mcsr/_0282_ ) );
AOI21_X1 \mcsr/_1770_ ( .A(\mcsr/_0761_ ), .B1(\mcsr/_0281_ ), .B2(\mcsr/_0282_ ), .ZN(\mcsr/_0072_ ) );
NAND2_X1 \mcsr/_1771_ ( .A1(\mcsr/_0764_ ), .A2(\mcsr/_0255_ ), .ZN(\mcsr/_0283_ ) );
NAND4_X1 \mcsr/_1772_ ( .A1(\mcsr/_0766_ ), .A2(\mcsr/_0897_ ), .A3(\mcsr/_0767_ ), .A4(\mcsr/_0768_ ), .ZN(\mcsr/_0284_ ) );
AOI21_X1 \mcsr/_1773_ ( .A(\mcsr/_0761_ ), .B1(\mcsr/_0283_ ), .B2(\mcsr/_0284_ ), .ZN(\mcsr/_0073_ ) );
NAND2_X1 \mcsr/_1774_ ( .A1(\mcsr/_0764_ ), .A2(\mcsr/_0225_ ), .ZN(\mcsr/_0285_ ) );
NAND4_X1 \mcsr/_1775_ ( .A1(\mcsr/_0766_ ), .A2(\mcsr/_0867_ ), .A3(\mcsr/_0767_ ), .A4(\mcsr/_0768_ ), .ZN(\mcsr/_0286_ ) );
AOI21_X1 \mcsr/_1776_ ( .A(\mcsr/_0761_ ), .B1(\mcsr/_0285_ ), .B2(\mcsr/_0286_ ), .ZN(\mcsr/_0074_ ) );
NAND2_X1 \mcsr/_1777_ ( .A1(\mcsr/_0764_ ), .A2(\mcsr/_0226_ ), .ZN(\mcsr/_0287_ ) );
NAND4_X1 \mcsr/_1778_ ( .A1(\mcsr/_0766_ ), .A2(\mcsr/_0868_ ), .A3(\mcsr/_0767_ ), .A4(\mcsr/_0768_ ), .ZN(\mcsr/_0288_ ) );
AOI21_X1 \mcsr/_1779_ ( .A(\mcsr/_0761_ ), .B1(\mcsr/_0287_ ), .B2(\mcsr/_0288_ ), .ZN(\mcsr/_0075_ ) );
NAND2_X1 \mcsr/_1780_ ( .A1(\mcsr/_0764_ ), .A2(\mcsr/_0227_ ), .ZN(\mcsr/_0289_ ) );
NAND4_X1 \mcsr/_1781_ ( .A1(\mcsr/_0766_ ), .A2(\mcsr/_0869_ ), .A3(\mcsr/_0767_ ), .A4(\mcsr/_0768_ ), .ZN(\mcsr/_0290_ ) );
AOI21_X1 \mcsr/_1782_ ( .A(\mcsr/_0761_ ), .B1(\mcsr/_0289_ ), .B2(\mcsr/_0290_ ), .ZN(\mcsr/_0076_ ) );
BUF_X4 \mcsr/_1783_ ( .A(\mcsr/_0679_ ), .Z(\mcsr/_0291_ ) );
BUF_X4 \mcsr/_1784_ ( .A(\mcsr/_0762_ ), .Z(\mcsr/_0292_ ) );
NAND2_X1 \mcsr/_1785_ ( .A1(\mcsr/_0292_ ), .A2(\mcsr/_0228_ ), .ZN(\mcsr/_0293_ ) );
BUF_X4 \mcsr/_1786_ ( .A(\mcsr/_0339_ ), .Z(\mcsr/_0294_ ) );
BUF_X4 \mcsr/_1787_ ( .A(\mcsr/_0341_ ), .Z(\mcsr/_0295_ ) );
BUF_X4 \mcsr/_1788_ ( .A(\mcsr/_0669_ ), .Z(\mcsr/_0296_ ) );
NAND4_X1 \mcsr/_1789_ ( .A1(\mcsr/_0294_ ), .A2(\mcsr/_0870_ ), .A3(\mcsr/_0295_ ), .A4(\mcsr/_0296_ ), .ZN(\mcsr/_0297_ ) );
AOI21_X1 \mcsr/_1790_ ( .A(\mcsr/_0291_ ), .B1(\mcsr/_0293_ ), .B2(\mcsr/_0297_ ), .ZN(\mcsr/_0077_ ) );
NAND2_X1 \mcsr/_1791_ ( .A1(\mcsr/_0292_ ), .A2(\mcsr/_0229_ ), .ZN(\mcsr/_0298_ ) );
NAND4_X1 \mcsr/_1792_ ( .A1(\mcsr/_0294_ ), .A2(\mcsr/_0871_ ), .A3(\mcsr/_0295_ ), .A4(\mcsr/_0296_ ), .ZN(\mcsr/_0299_ ) );
AOI21_X1 \mcsr/_1793_ ( .A(\mcsr/_0291_ ), .B1(\mcsr/_0298_ ), .B2(\mcsr/_0299_ ), .ZN(\mcsr/_0078_ ) );
NAND2_X1 \mcsr/_1794_ ( .A1(\mcsr/_0292_ ), .A2(\mcsr/_0230_ ), .ZN(\mcsr/_0300_ ) );
NAND4_X1 \mcsr/_1795_ ( .A1(\mcsr/_0294_ ), .A2(\mcsr/_0872_ ), .A3(\mcsr/_0295_ ), .A4(\mcsr/_0296_ ), .ZN(\mcsr/_0301_ ) );
AOI21_X1 \mcsr/_1796_ ( .A(\mcsr/_0291_ ), .B1(\mcsr/_0300_ ), .B2(\mcsr/_0301_ ), .ZN(\mcsr/_0079_ ) );
NAND2_X1 \mcsr/_1797_ ( .A1(\mcsr/_0292_ ), .A2(\mcsr/_0231_ ), .ZN(\mcsr/_0302_ ) );
NAND4_X1 \mcsr/_1798_ ( .A1(\mcsr/_0294_ ), .A2(\mcsr/_0873_ ), .A3(\mcsr/_0295_ ), .A4(\mcsr/_0296_ ), .ZN(\mcsr/_0303_ ) );
AOI21_X1 \mcsr/_1799_ ( .A(\mcsr/_0291_ ), .B1(\mcsr/_0302_ ), .B2(\mcsr/_0303_ ), .ZN(\mcsr/_0080_ ) );
NAND2_X1 \mcsr/_1800_ ( .A1(\mcsr/_0292_ ), .A2(\mcsr/_0232_ ), .ZN(\mcsr/_0304_ ) );
NAND4_X1 \mcsr/_1801_ ( .A1(\mcsr/_0294_ ), .A2(\mcsr/_0874_ ), .A3(\mcsr/_0295_ ), .A4(\mcsr/_0296_ ), .ZN(\mcsr/_0305_ ) );
AOI21_X1 \mcsr/_1802_ ( .A(\mcsr/_0291_ ), .B1(\mcsr/_0304_ ), .B2(\mcsr/_0305_ ), .ZN(\mcsr/_0081_ ) );
NAND2_X1 \mcsr/_1803_ ( .A1(\mcsr/_0292_ ), .A2(\mcsr/_0233_ ), .ZN(\mcsr/_0306_ ) );
NAND4_X1 \mcsr/_1804_ ( .A1(\mcsr/_0294_ ), .A2(\mcsr/_0875_ ), .A3(\mcsr/_0295_ ), .A4(\mcsr/_0296_ ), .ZN(\mcsr/_0307_ ) );
AOI21_X1 \mcsr/_1805_ ( .A(\mcsr/_0291_ ), .B1(\mcsr/_0306_ ), .B2(\mcsr/_0307_ ), .ZN(\mcsr/_0082_ ) );
NAND2_X1 \mcsr/_1806_ ( .A1(\mcsr/_0292_ ), .A2(\mcsr/_0234_ ), .ZN(\mcsr/_0308_ ) );
NAND4_X1 \mcsr/_1807_ ( .A1(\mcsr/_0294_ ), .A2(\mcsr/_0876_ ), .A3(\mcsr/_0295_ ), .A4(\mcsr/_0296_ ), .ZN(\mcsr/_0309_ ) );
AOI21_X1 \mcsr/_1808_ ( .A(\mcsr/_0291_ ), .B1(\mcsr/_0308_ ), .B2(\mcsr/_0309_ ), .ZN(\mcsr/_0083_ ) );
NAND2_X1 \mcsr/_1809_ ( .A1(\mcsr/_0292_ ), .A2(\mcsr/_0236_ ), .ZN(\mcsr/_0310_ ) );
NAND4_X1 \mcsr/_1810_ ( .A1(\mcsr/_0294_ ), .A2(\mcsr/_0878_ ), .A3(\mcsr/_0295_ ), .A4(\mcsr/_0296_ ), .ZN(\mcsr/_0311_ ) );
AOI21_X1 \mcsr/_1811_ ( .A(\mcsr/_0291_ ), .B1(\mcsr/_0310_ ), .B2(\mcsr/_0311_ ), .ZN(\mcsr/_0084_ ) );
NAND2_X1 \mcsr/_1812_ ( .A1(\mcsr/_0292_ ), .A2(\mcsr/_0237_ ), .ZN(\mcsr/_0312_ ) );
NAND4_X1 \mcsr/_1813_ ( .A1(\mcsr/_0294_ ), .A2(\mcsr/_0879_ ), .A3(\mcsr/_0295_ ), .A4(\mcsr/_0296_ ), .ZN(\mcsr/_0313_ ) );
AOI21_X1 \mcsr/_1814_ ( .A(\mcsr/_0291_ ), .B1(\mcsr/_0312_ ), .B2(\mcsr/_0313_ ), .ZN(\mcsr/_0085_ ) );
NAND2_X1 \mcsr/_1815_ ( .A1(\mcsr/_0292_ ), .A2(\mcsr/_0238_ ), .ZN(\mcsr/_0314_ ) );
NAND4_X1 \mcsr/_1816_ ( .A1(\mcsr/_0294_ ), .A2(\mcsr/_0880_ ), .A3(\mcsr/_0295_ ), .A4(\mcsr/_0296_ ), .ZN(\mcsr/_0315_ ) );
AOI21_X1 \mcsr/_1817_ ( .A(\mcsr/_0291_ ), .B1(\mcsr/_0314_ ), .B2(\mcsr/_0315_ ), .ZN(\mcsr/_0086_ ) );
NAND2_X1 \mcsr/_1818_ ( .A1(\mcsr/_0763_ ), .A2(\mcsr/_0239_ ), .ZN(\mcsr/_0316_ ) );
NAND4_X1 \mcsr/_1819_ ( .A1(\mcsr/_0754_ ), .A2(\mcsr/_0881_ ), .A3(\mcsr/_0755_ ), .A4(\mcsr/_0756_ ), .ZN(\mcsr/_0317_ ) );
AOI21_X1 \mcsr/_1820_ ( .A(\mcsr/_0760_ ), .B1(\mcsr/_0316_ ), .B2(\mcsr/_0317_ ), .ZN(\mcsr/_0087_ ) );
NAND2_X1 \mcsr/_1821_ ( .A1(\mcsr/_0763_ ), .A2(\mcsr/_0240_ ), .ZN(\mcsr/_0318_ ) );
NAND4_X1 \mcsr/_1822_ ( .A1(\mcsr/_0754_ ), .A2(\mcsr/_0882_ ), .A3(\mcsr/_0755_ ), .A4(\mcsr/_0756_ ), .ZN(\mcsr/_0319_ ) );
AOI21_X1 \mcsr/_1823_ ( .A(\mcsr/_0760_ ), .B1(\mcsr/_0318_ ), .B2(\mcsr/_0319_ ), .ZN(\mcsr/_0088_ ) );
NAND2_X1 \mcsr/_1824_ ( .A1(\mcsr/_0763_ ), .A2(\mcsr/_0241_ ), .ZN(\mcsr/_0320_ ) );
NAND4_X1 \mcsr/_1825_ ( .A1(\mcsr/_0754_ ), .A2(\mcsr/_0883_ ), .A3(\mcsr/_0755_ ), .A4(\mcsr/_0756_ ), .ZN(\mcsr/_0321_ ) );
AOI21_X1 \mcsr/_1826_ ( .A(\mcsr/_0760_ ), .B1(\mcsr/_0320_ ), .B2(\mcsr/_0321_ ), .ZN(\mcsr/_0089_ ) );
NAND2_X1 \mcsr/_1827_ ( .A1(\mcsr/_0763_ ), .A2(\mcsr/_0242_ ), .ZN(\mcsr/_0322_ ) );
NAND4_X1 \mcsr/_1828_ ( .A1(\mcsr/_0754_ ), .A2(\mcsr/_0884_ ), .A3(\mcsr/_0755_ ), .A4(\mcsr/_0756_ ), .ZN(\mcsr/_0323_ ) );
AOI21_X1 \mcsr/_1829_ ( .A(\mcsr/_0760_ ), .B1(\mcsr/_0322_ ), .B2(\mcsr/_0323_ ), .ZN(\mcsr/_0090_ ) );
NAND2_X1 \mcsr/_1830_ ( .A1(\mcsr/_0763_ ), .A2(\mcsr/_0243_ ), .ZN(\mcsr/_0324_ ) );
NAND4_X1 \mcsr/_1831_ ( .A1(\mcsr/_0754_ ), .A2(\mcsr/_0885_ ), .A3(\mcsr/_0755_ ), .A4(\mcsr/_0756_ ), .ZN(\mcsr/_0325_ ) );
AOI21_X1 \mcsr/_1832_ ( .A(\mcsr/_0760_ ), .B1(\mcsr/_0324_ ), .B2(\mcsr/_0325_ ), .ZN(\mcsr/_0091_ ) );
NAND2_X1 \mcsr/_1833_ ( .A1(\mcsr/_0763_ ), .A2(\mcsr/_0244_ ), .ZN(\mcsr/_0326_ ) );
NAND4_X1 \mcsr/_1834_ ( .A1(\mcsr/_0754_ ), .A2(\mcsr/_0886_ ), .A3(\mcsr/_0755_ ), .A4(\mcsr/_0756_ ), .ZN(\mcsr/_0327_ ) );
AOI21_X1 \mcsr/_1835_ ( .A(\mcsr/_0760_ ), .B1(\mcsr/_0326_ ), .B2(\mcsr/_0327_ ), .ZN(\mcsr/_0092_ ) );
NAND2_X1 \mcsr/_1836_ ( .A1(\mcsr/_0763_ ), .A2(\mcsr/_0245_ ), .ZN(\mcsr/_0328_ ) );
NAND4_X1 \mcsr/_1837_ ( .A1(\mcsr/_0754_ ), .A2(\mcsr/_0887_ ), .A3(\mcsr/_0755_ ), .A4(\mcsr/_0756_ ), .ZN(\mcsr/_0329_ ) );
AOI21_X1 \mcsr/_1838_ ( .A(\mcsr/_0760_ ), .B1(\mcsr/_0328_ ), .B2(\mcsr/_0329_ ), .ZN(\mcsr/_0093_ ) );
NAND2_X1 \mcsr/_1839_ ( .A1(\mcsr/_0763_ ), .A2(\mcsr/_0247_ ), .ZN(\mcsr/_0330_ ) );
NAND4_X1 \mcsr/_1840_ ( .A1(\mcsr/_0754_ ), .A2(\mcsr/_0889_ ), .A3(\mcsr/_0755_ ), .A4(\mcsr/_0756_ ), .ZN(\mcsr/_0331_ ) );
AOI21_X1 \mcsr/_1841_ ( .A(\mcsr/_0760_ ), .B1(\mcsr/_0330_ ), .B2(\mcsr/_0331_ ), .ZN(\mcsr/_0094_ ) );
NAND2_X1 \mcsr/_1842_ ( .A1(\mcsr/_0763_ ), .A2(\mcsr/_0248_ ), .ZN(\mcsr/_0332_ ) );
NAND4_X1 \mcsr/_1843_ ( .A1(\mcsr/_0754_ ), .A2(\mcsr/_0890_ ), .A3(\mcsr/_0755_ ), .A4(\mcsr/_0756_ ), .ZN(\mcsr/_0333_ ) );
AOI21_X1 \mcsr/_1844_ ( .A(\mcsr/_0760_ ), .B1(\mcsr/_0332_ ), .B2(\mcsr/_0333_ ), .ZN(\mcsr/_0095_ ) );
DFF_X1 \mcsr/_1845_ ( .CK(clk ), .D(\mcsr/_1027_ ), .Q(\mcsr/csr[1][0] ), .QN(\mcsr/_1026_ ) );
DFF_X1 \mcsr/_1846_ ( .CK(clk ), .D(\mcsr/_1028_ ), .Q(\mcsr/csr[1][1] ), .QN(\mcsr/_1025_ ) );
DFF_X1 \mcsr/_1847_ ( .CK(clk ), .D(\mcsr/_1029_ ), .Q(\mcsr/csr[1][2] ), .QN(\mcsr/_1024_ ) );
DFF_X1 \mcsr/_1848_ ( .CK(clk ), .D(\mcsr/_1030_ ), .Q(\mcsr/csr[1][3] ), .QN(\mcsr/_1023_ ) );
DFF_X1 \mcsr/_1849_ ( .CK(clk ), .D(\mcsr/_1031_ ), .Q(\mcsr/csr[1][4] ), .QN(\mcsr/_1022_ ) );
DFF_X1 \mcsr/_1850_ ( .CK(clk ), .D(\mcsr/_1032_ ), .Q(\mcsr/csr[1][5] ), .QN(\mcsr/_1021_ ) );
DFF_X1 \mcsr/_1851_ ( .CK(clk ), .D(\mcsr/_1033_ ), .Q(\mcsr/csr[1][6] ), .QN(\mcsr/_1020_ ) );
DFF_X1 \mcsr/_1852_ ( .CK(clk ), .D(\mcsr/_1034_ ), .Q(\mcsr/csr[1][7] ), .QN(\mcsr/_1019_ ) );
DFF_X1 \mcsr/_1853_ ( .CK(clk ), .D(\mcsr/_1035_ ), .Q(\mcsr/csr[1][8] ), .QN(\mcsr/_1018_ ) );
DFF_X1 \mcsr/_1854_ ( .CK(clk ), .D(\mcsr/_1036_ ), .Q(\mcsr/csr[1][9] ), .QN(\mcsr/_1017_ ) );
DFF_X1 \mcsr/_1855_ ( .CK(clk ), .D(\mcsr/_1037_ ), .Q(\mcsr/csr[1][10] ), .QN(\mcsr/_1016_ ) );
DFF_X1 \mcsr/_1856_ ( .CK(clk ), .D(\mcsr/_1038_ ), .Q(\mcsr/csr[1][11] ), .QN(\mcsr/_1015_ ) );
DFF_X1 \mcsr/_1857_ ( .CK(clk ), .D(\mcsr/_1039_ ), .Q(\mcsr/csr[1][12] ), .QN(\mcsr/_1014_ ) );
DFF_X1 \mcsr/_1858_ ( .CK(clk ), .D(\mcsr/_1040_ ), .Q(\mcsr/csr[1][13] ), .QN(\mcsr/_1013_ ) );
DFF_X1 \mcsr/_1859_ ( .CK(clk ), .D(\mcsr/_1041_ ), .Q(\mcsr/csr[1][14] ), .QN(\mcsr/_1012_ ) );
DFF_X1 \mcsr/_1860_ ( .CK(clk ), .D(\mcsr/_1042_ ), .Q(\mcsr/csr[1][15] ), .QN(\mcsr/_1011_ ) );
DFF_X1 \mcsr/_1861_ ( .CK(clk ), .D(\mcsr/_1043_ ), .Q(\mcsr/csr[1][16] ), .QN(\mcsr/_1010_ ) );
DFF_X1 \mcsr/_1862_ ( .CK(clk ), .D(\mcsr/_1044_ ), .Q(\mcsr/csr[1][17] ), .QN(\mcsr/_1009_ ) );
DFF_X1 \mcsr/_1863_ ( .CK(clk ), .D(\mcsr/_1045_ ), .Q(\mcsr/csr[1][18] ), .QN(\mcsr/_1008_ ) );
DFF_X1 \mcsr/_1864_ ( .CK(clk ), .D(\mcsr/_1046_ ), .Q(\mcsr/csr[1][19] ), .QN(\mcsr/_1007_ ) );
DFF_X1 \mcsr/_1865_ ( .CK(clk ), .D(\mcsr/_1047_ ), .Q(\mcsr/csr[1][20] ), .QN(\mcsr/_1006_ ) );
DFF_X1 \mcsr/_1866_ ( .CK(clk ), .D(\mcsr/_1048_ ), .Q(\mcsr/csr[1][21] ), .QN(\mcsr/_1005_ ) );
DFF_X1 \mcsr/_1867_ ( .CK(clk ), .D(\mcsr/_1049_ ), .Q(\mcsr/csr[1][22] ), .QN(\mcsr/_1004_ ) );
DFF_X1 \mcsr/_1868_ ( .CK(clk ), .D(\mcsr/_1050_ ), .Q(\mcsr/csr[1][23] ), .QN(\mcsr/_1003_ ) );
DFF_X1 \mcsr/_1869_ ( .CK(clk ), .D(\mcsr/_1051_ ), .Q(\mcsr/csr[1][24] ), .QN(\mcsr/_1002_ ) );
DFF_X1 \mcsr/_1870_ ( .CK(clk ), .D(\mcsr/_1052_ ), .Q(\mcsr/csr[1][25] ), .QN(\mcsr/_1001_ ) );
DFF_X1 \mcsr/_1871_ ( .CK(clk ), .D(\mcsr/_1053_ ), .Q(\mcsr/csr[1][26] ), .QN(\mcsr/_1000_ ) );
DFF_X1 \mcsr/_1872_ ( .CK(clk ), .D(\mcsr/_1054_ ), .Q(\mcsr/csr[1][27] ), .QN(\mcsr/_0999_ ) );
DFF_X1 \mcsr/_1873_ ( .CK(clk ), .D(\mcsr/_1055_ ), .Q(\mcsr/csr[1][28] ), .QN(\mcsr/_0998_ ) );
DFF_X1 \mcsr/_1874_ ( .CK(clk ), .D(\mcsr/_1056_ ), .Q(\mcsr/csr[1][29] ), .QN(\mcsr/_0997_ ) );
DFF_X1 \mcsr/_1875_ ( .CK(clk ), .D(\mcsr/_1057_ ), .Q(\mcsr/csr[1][30] ), .QN(\mcsr/_0996_ ) );
DFF_X1 \mcsr/_1876_ ( .CK(clk ), .D(\mcsr/_1058_ ), .Q(\mcsr/csr[1][31] ), .QN(\mcsr/_0995_ ) );
DFF_X1 \mcsr/_1877_ ( .CK(clk ), .D(\mcsr/_1059_ ), .Q(\mcsr/csr[2][0] ), .QN(\mcsr/_0994_ ) );
DFF_X1 \mcsr/_1878_ ( .CK(clk ), .D(\mcsr/_1060_ ), .Q(\mcsr/csr[2][1] ), .QN(\mcsr/_0993_ ) );
DFF_X1 \mcsr/_1879_ ( .CK(clk ), .D(\mcsr/_1061_ ), .Q(\mcsr/csr[2][2] ), .QN(\mcsr/_0992_ ) );
DFF_X1 \mcsr/_1880_ ( .CK(clk ), .D(\mcsr/_1062_ ), .Q(\mcsr/csr[2][3] ), .QN(\mcsr/_0991_ ) );
DFF_X1 \mcsr/_1881_ ( .CK(clk ), .D(\mcsr/_1063_ ), .Q(\mcsr/csr[2][4] ), .QN(\mcsr/_0990_ ) );
DFF_X1 \mcsr/_1882_ ( .CK(clk ), .D(\mcsr/_1064_ ), .Q(\mcsr/csr[2][5] ), .QN(\mcsr/_0989_ ) );
DFF_X1 \mcsr/_1883_ ( .CK(clk ), .D(\mcsr/_1065_ ), .Q(\mcsr/csr[2][6] ), .QN(\mcsr/_0988_ ) );
DFF_X1 \mcsr/_1884_ ( .CK(clk ), .D(\mcsr/_1066_ ), .Q(\mcsr/csr[2][7] ), .QN(\mcsr/_0987_ ) );
DFF_X1 \mcsr/_1885_ ( .CK(clk ), .D(\mcsr/_1067_ ), .Q(\mcsr/csr[2][8] ), .QN(\mcsr/_0986_ ) );
DFF_X1 \mcsr/_1886_ ( .CK(clk ), .D(\mcsr/_1068_ ), .Q(\mcsr/csr[2][9] ), .QN(\mcsr/_0985_ ) );
DFF_X1 \mcsr/_1887_ ( .CK(clk ), .D(\mcsr/_1069_ ), .Q(\mcsr/csr[2][10] ), .QN(\mcsr/_0984_ ) );
DFF_X1 \mcsr/_1888_ ( .CK(clk ), .D(\mcsr/_1070_ ), .Q(\mcsr/csr[2][11] ), .QN(\mcsr/_0983_ ) );
DFF_X1 \mcsr/_1889_ ( .CK(clk ), .D(\mcsr/_1071_ ), .Q(\mcsr/csr[2][12] ), .QN(\mcsr/_0982_ ) );
DFF_X1 \mcsr/_1890_ ( .CK(clk ), .D(\mcsr/_1072_ ), .Q(\mcsr/csr[2][13] ), .QN(\mcsr/_0981_ ) );
DFF_X1 \mcsr/_1891_ ( .CK(clk ), .D(\mcsr/_1073_ ), .Q(\mcsr/csr[2][14] ), .QN(\mcsr/_0980_ ) );
DFF_X1 \mcsr/_1892_ ( .CK(clk ), .D(\mcsr/_1074_ ), .Q(\mcsr/csr[2][15] ), .QN(\mcsr/_0979_ ) );
DFF_X1 \mcsr/_1893_ ( .CK(clk ), .D(\mcsr/_1075_ ), .Q(\mcsr/csr[2][16] ), .QN(\mcsr/_0978_ ) );
DFF_X1 \mcsr/_1894_ ( .CK(clk ), .D(\mcsr/_1076_ ), .Q(\mcsr/csr[2][17] ), .QN(\mcsr/_0977_ ) );
DFF_X1 \mcsr/_1895_ ( .CK(clk ), .D(\mcsr/_1077_ ), .Q(\mcsr/csr[2][18] ), .QN(\mcsr/_0976_ ) );
DFF_X1 \mcsr/_1896_ ( .CK(clk ), .D(\mcsr/_1078_ ), .Q(\mcsr/csr[2][19] ), .QN(\mcsr/_0975_ ) );
DFF_X1 \mcsr/_1897_ ( .CK(clk ), .D(\mcsr/_1079_ ), .Q(\mcsr/csr[2][20] ), .QN(\mcsr/_0974_ ) );
DFF_X1 \mcsr/_1898_ ( .CK(clk ), .D(\mcsr/_1080_ ), .Q(\mcsr/csr[2][21] ), .QN(\mcsr/_0973_ ) );
DFF_X1 \mcsr/_1899_ ( .CK(clk ), .D(\mcsr/_1081_ ), .Q(\mcsr/csr[2][22] ), .QN(\mcsr/_0972_ ) );
DFF_X1 \mcsr/_1900_ ( .CK(clk ), .D(\mcsr/_1082_ ), .Q(\mcsr/csr[2][23] ), .QN(\mcsr/_0971_ ) );
DFF_X1 \mcsr/_1901_ ( .CK(clk ), .D(\mcsr/_1083_ ), .Q(\mcsr/csr[2][24] ), .QN(\mcsr/_0970_ ) );
DFF_X1 \mcsr/_1902_ ( .CK(clk ), .D(\mcsr/_1084_ ), .Q(\mcsr/csr[2][25] ), .QN(\mcsr/_0969_ ) );
DFF_X1 \mcsr/_1903_ ( .CK(clk ), .D(\mcsr/_1085_ ), .Q(\mcsr/csr[2][26] ), .QN(\mcsr/_0968_ ) );
DFF_X1 \mcsr/_1904_ ( .CK(clk ), .D(\mcsr/_1086_ ), .Q(\mcsr/csr[2][27] ), .QN(\mcsr/_0967_ ) );
DFF_X1 \mcsr/_1905_ ( .CK(clk ), .D(\mcsr/_1087_ ), .Q(\mcsr/csr[2][28] ), .QN(\mcsr/_0966_ ) );
DFF_X1 \mcsr/_1906_ ( .CK(clk ), .D(\mcsr/_1088_ ), .Q(\mcsr/csr[2][29] ), .QN(\mcsr/_0965_ ) );
DFF_X1 \mcsr/_1907_ ( .CK(clk ), .D(\mcsr/_1089_ ), .Q(\mcsr/csr[2][30] ), .QN(\mcsr/_0964_ ) );
DFF_X1 \mcsr/_1908_ ( .CK(clk ), .D(\mcsr/_1090_ ), .Q(\mcsr/csr[2][31] ), .QN(\mcsr/_0963_ ) );
DFF_X1 \mcsr/_1909_ ( .CK(clk ), .D(\mcsr/_1091_ ), .Q(\mcsr/csr[3][0] ), .QN(\mcsr/_0962_ ) );
DFF_X1 \mcsr/_1910_ ( .CK(clk ), .D(\mcsr/_1092_ ), .Q(\mcsr/csr[3][1] ), .QN(\mcsr/_0961_ ) );
DFF_X1 \mcsr/_1911_ ( .CK(clk ), .D(\mcsr/_1093_ ), .Q(\mcsr/csr[3][2] ), .QN(\mcsr/_0960_ ) );
DFF_X1 \mcsr/_1912_ ( .CK(clk ), .D(\mcsr/_1094_ ), .Q(\mcsr/csr[3][3] ), .QN(\mcsr/_0959_ ) );
DFF_X1 \mcsr/_1913_ ( .CK(clk ), .D(\mcsr/_1095_ ), .Q(\mcsr/csr[3][4] ), .QN(\mcsr/_0958_ ) );
DFF_X1 \mcsr/_1914_ ( .CK(clk ), .D(\mcsr/_1096_ ), .Q(\mcsr/csr[3][5] ), .QN(\mcsr/_0957_ ) );
DFF_X1 \mcsr/_1915_ ( .CK(clk ), .D(\mcsr/_1097_ ), .Q(\mcsr/csr[3][6] ), .QN(\mcsr/_0956_ ) );
DFF_X1 \mcsr/_1916_ ( .CK(clk ), .D(\mcsr/_1098_ ), .Q(\mcsr/csr[3][7] ), .QN(\mcsr/_0955_ ) );
DFF_X1 \mcsr/_1917_ ( .CK(clk ), .D(\mcsr/_1099_ ), .Q(\mcsr/csr[3][8] ), .QN(\mcsr/_0954_ ) );
DFF_X1 \mcsr/_1918_ ( .CK(clk ), .D(\mcsr/_1100_ ), .Q(\mcsr/csr[3][9] ), .QN(\mcsr/_0953_ ) );
DFF_X1 \mcsr/_1919_ ( .CK(clk ), .D(\mcsr/_1101_ ), .Q(\mcsr/csr[3][10] ), .QN(\mcsr/_0952_ ) );
DFF_X1 \mcsr/_1920_ ( .CK(clk ), .D(\mcsr/_1102_ ), .Q(\mcsr/csr[3][11] ), .QN(\mcsr/_0951_ ) );
DFF_X1 \mcsr/_1921_ ( .CK(clk ), .D(\mcsr/_1103_ ), .Q(\mcsr/csr[3][12] ), .QN(\mcsr/_0950_ ) );
DFF_X1 \mcsr/_1922_ ( .CK(clk ), .D(\mcsr/_1104_ ), .Q(\mcsr/csr[3][13] ), .QN(\mcsr/_0949_ ) );
DFF_X1 \mcsr/_1923_ ( .CK(clk ), .D(\mcsr/_1105_ ), .Q(\mcsr/csr[3][14] ), .QN(\mcsr/_0948_ ) );
DFF_X1 \mcsr/_1924_ ( .CK(clk ), .D(\mcsr/_1106_ ), .Q(\mcsr/csr[3][15] ), .QN(\mcsr/_0947_ ) );
DFF_X1 \mcsr/_1925_ ( .CK(clk ), .D(\mcsr/_1107_ ), .Q(\mcsr/csr[3][16] ), .QN(\mcsr/_0946_ ) );
DFF_X1 \mcsr/_1926_ ( .CK(clk ), .D(\mcsr/_1108_ ), .Q(\mcsr/csr[3][17] ), .QN(\mcsr/_0945_ ) );
DFF_X1 \mcsr/_1927_ ( .CK(clk ), .D(\mcsr/_1109_ ), .Q(\mcsr/csr[3][18] ), .QN(\mcsr/_0944_ ) );
DFF_X1 \mcsr/_1928_ ( .CK(clk ), .D(\mcsr/_1110_ ), .Q(\mcsr/csr[3][19] ), .QN(\mcsr/_0943_ ) );
DFF_X1 \mcsr/_1929_ ( .CK(clk ), .D(\mcsr/_1111_ ), .Q(\mcsr/csr[3][20] ), .QN(\mcsr/_0942_ ) );
DFF_X1 \mcsr/_1930_ ( .CK(clk ), .D(\mcsr/_1112_ ), .Q(\mcsr/csr[3][21] ), .QN(\mcsr/_0941_ ) );
DFF_X1 \mcsr/_1931_ ( .CK(clk ), .D(\mcsr/_1113_ ), .Q(\mcsr/csr[3][22] ), .QN(\mcsr/_0940_ ) );
DFF_X1 \mcsr/_1932_ ( .CK(clk ), .D(\mcsr/_1114_ ), .Q(\mcsr/csr[3][23] ), .QN(\mcsr/_0939_ ) );
DFF_X1 \mcsr/_1933_ ( .CK(clk ), .D(\mcsr/_1115_ ), .Q(\mcsr/csr[3][24] ), .QN(\mcsr/_0938_ ) );
DFF_X1 \mcsr/_1934_ ( .CK(clk ), .D(\mcsr/_1116_ ), .Q(\mcsr/csr[3][25] ), .QN(\mcsr/_0937_ ) );
DFF_X1 \mcsr/_1935_ ( .CK(clk ), .D(\mcsr/_1117_ ), .Q(\mcsr/csr[3][26] ), .QN(\mcsr/_0936_ ) );
DFF_X1 \mcsr/_1936_ ( .CK(clk ), .D(\mcsr/_1118_ ), .Q(\mcsr/csr[3][27] ), .QN(\mcsr/_0935_ ) );
DFF_X1 \mcsr/_1937_ ( .CK(clk ), .D(\mcsr/_1119_ ), .Q(\mcsr/csr[3][28] ), .QN(\mcsr/_0934_ ) );
DFF_X1 \mcsr/_1938_ ( .CK(clk ), .D(\mcsr/_1120_ ), .Q(\mcsr/csr[3][29] ), .QN(\mcsr/_0933_ ) );
DFF_X1 \mcsr/_1939_ ( .CK(clk ), .D(\mcsr/_1121_ ), .Q(\mcsr/csr[3][30] ), .QN(\mcsr/_0932_ ) );
DFF_X1 \mcsr/_1940_ ( .CK(clk ), .D(\mcsr/_1122_ ), .Q(\mcsr/csr[3][31] ), .QN(\mcsr/_0931_ ) );
DFF_X1 \mcsr/_1941_ ( .CK(clk ), .D(\mcsr/_1123_ ), .Q(\mcsr/csr[0][0] ), .QN(\mcsr/_0930_ ) );
DFF_X1 \mcsr/_1942_ ( .CK(clk ), .D(\mcsr/_1124_ ), .Q(\mcsr/csr[0][1] ), .QN(\mcsr/_0929_ ) );
DFF_X1 \mcsr/_1943_ ( .CK(clk ), .D(\mcsr/_1125_ ), .Q(\mcsr/csr[0][2] ), .QN(\mcsr/_0928_ ) );
DFF_X1 \mcsr/_1944_ ( .CK(clk ), .D(\mcsr/_1126_ ), .Q(\mcsr/csr[0][3] ), .QN(\mcsr/_0927_ ) );
DFF_X1 \mcsr/_1945_ ( .CK(clk ), .D(\mcsr/_1127_ ), .Q(\mcsr/csr[0][4] ), .QN(\mcsr/_0926_ ) );
DFF_X1 \mcsr/_1946_ ( .CK(clk ), .D(\mcsr/_1128_ ), .Q(\mcsr/csr[0][5] ), .QN(\mcsr/_0925_ ) );
DFF_X1 \mcsr/_1947_ ( .CK(clk ), .D(\mcsr/_1129_ ), .Q(\mcsr/csr[0][6] ), .QN(\mcsr/_0924_ ) );
DFF_X1 \mcsr/_1948_ ( .CK(clk ), .D(\mcsr/_1130_ ), .Q(\mcsr/csr[0][7] ), .QN(\mcsr/_0923_ ) );
DFF_X1 \mcsr/_1949_ ( .CK(clk ), .D(\mcsr/_1131_ ), .Q(\mcsr/csr[0][8] ), .QN(\mcsr/_0922_ ) );
DFF_X1 \mcsr/_1950_ ( .CK(clk ), .D(\mcsr/_1132_ ), .Q(\mcsr/csr[0][9] ), .QN(\mcsr/_0921_ ) );
DFF_X1 \mcsr/_1951_ ( .CK(clk ), .D(\mcsr/_1133_ ), .Q(\mcsr/csr[0][10] ), .QN(\mcsr/_0920_ ) );
DFF_X1 \mcsr/_1952_ ( .CK(clk ), .D(\mcsr/_1134_ ), .Q(\mcsr/csr[0][11] ), .QN(\mcsr/_0919_ ) );
DFF_X1 \mcsr/_1953_ ( .CK(clk ), .D(\mcsr/_1135_ ), .Q(\mcsr/csr[0][12] ), .QN(\mcsr/_0918_ ) );
DFF_X1 \mcsr/_1954_ ( .CK(clk ), .D(\mcsr/_1136_ ), .Q(\mcsr/csr[0][13] ), .QN(\mcsr/_0917_ ) );
DFF_X1 \mcsr/_1955_ ( .CK(clk ), .D(\mcsr/_1137_ ), .Q(\mcsr/csr[0][14] ), .QN(\mcsr/_0916_ ) );
DFF_X1 \mcsr/_1956_ ( .CK(clk ), .D(\mcsr/_1138_ ), .Q(\mcsr/csr[0][15] ), .QN(\mcsr/_0915_ ) );
DFF_X1 \mcsr/_1957_ ( .CK(clk ), .D(\mcsr/_1139_ ), .Q(\mcsr/csr[0][16] ), .QN(\mcsr/_0914_ ) );
DFF_X1 \mcsr/_1958_ ( .CK(clk ), .D(\mcsr/_1140_ ), .Q(\mcsr/csr[0][17] ), .QN(\mcsr/_0913_ ) );
DFF_X1 \mcsr/_1959_ ( .CK(clk ), .D(\mcsr/_1141_ ), .Q(\mcsr/csr[0][18] ), .QN(\mcsr/_0912_ ) );
DFF_X1 \mcsr/_1960_ ( .CK(clk ), .D(\mcsr/_1142_ ), .Q(\mcsr/csr[0][19] ), .QN(\mcsr/_0911_ ) );
DFF_X1 \mcsr/_1961_ ( .CK(clk ), .D(\mcsr/_1143_ ), .Q(\mcsr/csr[0][20] ), .QN(\mcsr/_0910_ ) );
DFF_X1 \mcsr/_1962_ ( .CK(clk ), .D(\mcsr/_1144_ ), .Q(\mcsr/csr[0][21] ), .QN(\mcsr/_0909_ ) );
DFF_X1 \mcsr/_1963_ ( .CK(clk ), .D(\mcsr/_1145_ ), .Q(\mcsr/csr[0][22] ), .QN(\mcsr/_0908_ ) );
DFF_X1 \mcsr/_1964_ ( .CK(clk ), .D(\mcsr/_1146_ ), .Q(\mcsr/csr[0][23] ), .QN(\mcsr/_0907_ ) );
DFF_X1 \mcsr/_1965_ ( .CK(clk ), .D(\mcsr/_1147_ ), .Q(\mcsr/csr[0][24] ), .QN(\mcsr/_0906_ ) );
DFF_X1 \mcsr/_1966_ ( .CK(clk ), .D(\mcsr/_1148_ ), .Q(\mcsr/csr[0][25] ), .QN(\mcsr/_0905_ ) );
DFF_X1 \mcsr/_1967_ ( .CK(clk ), .D(\mcsr/_1149_ ), .Q(\mcsr/csr[0][26] ), .QN(\mcsr/_0904_ ) );
DFF_X1 \mcsr/_1968_ ( .CK(clk ), .D(\mcsr/_1150_ ), .Q(\mcsr/csr[0][27] ), .QN(\mcsr/_0903_ ) );
DFF_X1 \mcsr/_1969_ ( .CK(clk ), .D(\mcsr/_1151_ ), .Q(\mcsr/csr[0][28] ), .QN(\mcsr/_0902_ ) );
DFF_X1 \mcsr/_1970_ ( .CK(clk ), .D(\mcsr/_1152_ ), .Q(\mcsr/csr[0][29] ), .QN(\mcsr/_0901_ ) );
DFF_X1 \mcsr/_1971_ ( .CK(clk ), .D(\mcsr/_1153_ ), .Q(\mcsr/csr[0][30] ), .QN(\mcsr/_0900_ ) );
DFF_X1 \mcsr/_1972_ ( .CK(clk ), .D(\mcsr/_1154_ ), .Q(\mcsr/csr[0][31] ), .QN(\mcsr/_0899_ ) );
BUF_X1 \mcsr/_1973_ ( .A(csr_wen ), .Z(\mcsr/_0898_ ) );
BUF_X1 \mcsr/_1974_ ( .A(lsu_finish ), .Z(\mcsr/_0271_ ) );
BUF_X1 \mcsr/_1975_ ( .A(\csr_ctl[0] ), .Z(\mcsr/_0268_ ) );
BUF_X1 \mcsr/_1976_ ( .A(\csr_ctl[1] ), .Z(\mcsr/_0269_ ) );
BUF_X1 \mcsr/_1977_ ( .A(\csr_ctl[2] ), .Z(\mcsr/_0270_ ) );
BUF_X1 \mcsr/_1978_ ( .A(\imm[1] ), .Z(\mcsr/_0259_ ) );
BUF_X1 \mcsr/_1979_ ( .A(\imm[0] ), .Z(\mcsr/_0256_ ) );
BUF_X1 \mcsr/_1980_ ( .A(\imm[3] ), .Z(\mcsr/_0261_ ) );
BUF_X1 \mcsr/_1981_ ( .A(\imm[2] ), .Z(\mcsr/_0260_ ) );
BUF_X1 \mcsr/_1982_ ( .A(\imm[5] ), .Z(\mcsr/_0263_ ) );
BUF_X1 \mcsr/_1983_ ( .A(\imm[4] ), .Z(\mcsr/_0262_ ) );
BUF_X1 \mcsr/_1984_ ( .A(\imm[7] ), .Z(\mcsr/_0265_ ) );
BUF_X1 \mcsr/_1985_ ( .A(\imm[6] ), .Z(\mcsr/_0264_ ) );
BUF_X1 \mcsr/_1986_ ( .A(\imm[9] ), .Z(\mcsr/_0267_ ) );
BUF_X1 \mcsr/_1987_ ( .A(\imm[8] ), .Z(\mcsr/_0266_ ) );
BUF_X1 \mcsr/_1988_ ( .A(\imm[11] ), .Z(\mcsr/_0258_ ) );
BUF_X1 \mcsr/_1989_ ( .A(\imm[10] ), .Z(\mcsr/_0257_ ) );
BUF_X1 \mcsr/_1990_ ( .A(\mcsr/csr[1][0] ), .Z(\mcsr/_0160_ ) );
BUF_X1 \mcsr/_1991_ ( .A(\mcsr/csr[0][0] ), .Z(\mcsr/_0128_ ) );
BUF_X1 \mcsr/_1992_ ( .A(\mcsr/csr[3][0] ), .Z(\mcsr/_0224_ ) );
BUF_X1 \mcsr/_1993_ ( .A(\mcsr/csr[2][0] ), .Z(\mcsr/_0192_ ) );
BUF_X1 \mcsr/_1994_ ( .A(\mcsr/_0802_ ), .Z(\csr_rdata[0] ) );
BUF_X1 \mcsr/_1995_ ( .A(\mcsr/csr[1][1] ), .Z(\mcsr/_0171_ ) );
BUF_X1 \mcsr/_1996_ ( .A(\mcsr/csr[0][1] ), .Z(\mcsr/_0139_ ) );
BUF_X1 \mcsr/_1997_ ( .A(\mcsr/csr[3][1] ), .Z(\mcsr/_0235_ ) );
BUF_X1 \mcsr/_1998_ ( .A(\mcsr/csr[2][1] ), .Z(\mcsr/_0203_ ) );
BUF_X1 \mcsr/_1999_ ( .A(\mcsr/_0813_ ), .Z(\csr_rdata[1] ) );
BUF_X1 \mcsr/_2000_ ( .A(\mcsr/csr[1][2] ), .Z(\mcsr/_0182_ ) );
BUF_X1 \mcsr/_2001_ ( .A(\mcsr/csr[0][2] ), .Z(\mcsr/_0150_ ) );
BUF_X1 \mcsr/_2002_ ( .A(\mcsr/csr[3][2] ), .Z(\mcsr/_0246_ ) );
BUF_X1 \mcsr/_2003_ ( .A(\mcsr/csr[2][2] ), .Z(\mcsr/_0214_ ) );
BUF_X1 \mcsr/_2004_ ( .A(\mcsr/_0824_ ), .Z(\csr_rdata[2] ) );
BUF_X1 \mcsr/_2005_ ( .A(\mcsr/csr[1][3] ), .Z(\mcsr/_0185_ ) );
BUF_X1 \mcsr/_2006_ ( .A(\mcsr/csr[0][3] ), .Z(\mcsr/_0153_ ) );
BUF_X1 \mcsr/_2007_ ( .A(\mcsr/csr[3][3] ), .Z(\mcsr/_0249_ ) );
BUF_X1 \mcsr/_2008_ ( .A(\mcsr/csr[2][3] ), .Z(\mcsr/_0217_ ) );
BUF_X1 \mcsr/_2009_ ( .A(\mcsr/_0827_ ), .Z(\csr_rdata[3] ) );
BUF_X1 \mcsr/_2010_ ( .A(\mcsr/csr[1][4] ), .Z(\mcsr/_0186_ ) );
BUF_X1 \mcsr/_2011_ ( .A(\mcsr/csr[0][4] ), .Z(\mcsr/_0154_ ) );
BUF_X1 \mcsr/_2012_ ( .A(\mcsr/csr[3][4] ), .Z(\mcsr/_0250_ ) );
BUF_X1 \mcsr/_2013_ ( .A(\mcsr/csr[2][4] ), .Z(\mcsr/_0218_ ) );
BUF_X1 \mcsr/_2014_ ( .A(\mcsr/_0828_ ), .Z(\csr_rdata[4] ) );
BUF_X1 \mcsr/_2015_ ( .A(\mcsr/csr[1][5] ), .Z(\mcsr/_0187_ ) );
BUF_X1 \mcsr/_2016_ ( .A(\mcsr/csr[0][5] ), .Z(\mcsr/_0155_ ) );
BUF_X1 \mcsr/_2017_ ( .A(\mcsr/csr[3][5] ), .Z(\mcsr/_0251_ ) );
BUF_X1 \mcsr/_2018_ ( .A(\mcsr/csr[2][5] ), .Z(\mcsr/_0219_ ) );
BUF_X1 \mcsr/_2019_ ( .A(\mcsr/_0829_ ), .Z(\csr_rdata[5] ) );
BUF_X1 \mcsr/_2020_ ( .A(\mcsr/csr[1][6] ), .Z(\mcsr/_0188_ ) );
BUF_X1 \mcsr/_2021_ ( .A(\mcsr/csr[0][6] ), .Z(\mcsr/_0156_ ) );
BUF_X1 \mcsr/_2022_ ( .A(\mcsr/csr[3][6] ), .Z(\mcsr/_0252_ ) );
BUF_X1 \mcsr/_2023_ ( .A(\mcsr/csr[2][6] ), .Z(\mcsr/_0220_ ) );
BUF_X1 \mcsr/_2024_ ( .A(\mcsr/_0830_ ), .Z(\csr_rdata[6] ) );
BUF_X1 \mcsr/_2025_ ( .A(\mcsr/csr[1][7] ), .Z(\mcsr/_0189_ ) );
BUF_X1 \mcsr/_2026_ ( .A(\mcsr/csr[0][7] ), .Z(\mcsr/_0157_ ) );
BUF_X1 \mcsr/_2027_ ( .A(\mcsr/csr[3][7] ), .Z(\mcsr/_0253_ ) );
BUF_X1 \mcsr/_2028_ ( .A(\mcsr/csr[2][7] ), .Z(\mcsr/_0221_ ) );
BUF_X1 \mcsr/_2029_ ( .A(\mcsr/_0831_ ), .Z(\csr_rdata[7] ) );
BUF_X1 \mcsr/_2030_ ( .A(\mcsr/csr[1][8] ), .Z(\mcsr/_0190_ ) );
BUF_X1 \mcsr/_2031_ ( .A(\mcsr/csr[0][8] ), .Z(\mcsr/_0158_ ) );
BUF_X1 \mcsr/_2032_ ( .A(\mcsr/csr[3][8] ), .Z(\mcsr/_0254_ ) );
BUF_X1 \mcsr/_2033_ ( .A(\mcsr/csr[2][8] ), .Z(\mcsr/_0222_ ) );
BUF_X1 \mcsr/_2034_ ( .A(\mcsr/_0832_ ), .Z(\csr_rdata[8] ) );
BUF_X1 \mcsr/_2035_ ( .A(\mcsr/csr[1][9] ), .Z(\mcsr/_0191_ ) );
BUF_X1 \mcsr/_2036_ ( .A(\mcsr/csr[0][9] ), .Z(\mcsr/_0159_ ) );
BUF_X1 \mcsr/_2037_ ( .A(\mcsr/csr[3][9] ), .Z(\mcsr/_0255_ ) );
BUF_X1 \mcsr/_2038_ ( .A(\mcsr/csr[2][9] ), .Z(\mcsr/_0223_ ) );
BUF_X1 \mcsr/_2039_ ( .A(\mcsr/_0833_ ), .Z(\csr_rdata[9] ) );
BUF_X1 \mcsr/_2040_ ( .A(\mcsr/csr[1][10] ), .Z(\mcsr/_0161_ ) );
BUF_X1 \mcsr/_2041_ ( .A(\mcsr/csr[0][10] ), .Z(\mcsr/_0129_ ) );
BUF_X1 \mcsr/_2042_ ( .A(\mcsr/csr[3][10] ), .Z(\mcsr/_0225_ ) );
BUF_X1 \mcsr/_2043_ ( .A(\mcsr/csr[2][10] ), .Z(\mcsr/_0193_ ) );
BUF_X1 \mcsr/_2044_ ( .A(\mcsr/_0803_ ), .Z(\csr_rdata[10] ) );
BUF_X1 \mcsr/_2045_ ( .A(\mcsr/csr[1][11] ), .Z(\mcsr/_0162_ ) );
BUF_X1 \mcsr/_2046_ ( .A(\mcsr/csr[0][11] ), .Z(\mcsr/_0130_ ) );
BUF_X1 \mcsr/_2047_ ( .A(\mcsr/csr[3][11] ), .Z(\mcsr/_0226_ ) );
BUF_X1 \mcsr/_2048_ ( .A(\mcsr/csr[2][11] ), .Z(\mcsr/_0194_ ) );
BUF_X1 \mcsr/_2049_ ( .A(\mcsr/_0804_ ), .Z(\csr_rdata[11] ) );
BUF_X1 \mcsr/_2050_ ( .A(\mcsr/csr[1][12] ), .Z(\mcsr/_0163_ ) );
BUF_X1 \mcsr/_2051_ ( .A(\mcsr/csr[0][12] ), .Z(\mcsr/_0131_ ) );
BUF_X1 \mcsr/_2052_ ( .A(\mcsr/csr[3][12] ), .Z(\mcsr/_0227_ ) );
BUF_X1 \mcsr/_2053_ ( .A(\mcsr/csr[2][12] ), .Z(\mcsr/_0195_ ) );
BUF_X1 \mcsr/_2054_ ( .A(\mcsr/_0805_ ), .Z(\csr_rdata[12] ) );
BUF_X1 \mcsr/_2055_ ( .A(\mcsr/csr[1][13] ), .Z(\mcsr/_0164_ ) );
BUF_X1 \mcsr/_2056_ ( .A(\mcsr/csr[0][13] ), .Z(\mcsr/_0132_ ) );
BUF_X1 \mcsr/_2057_ ( .A(\mcsr/csr[3][13] ), .Z(\mcsr/_0228_ ) );
BUF_X1 \mcsr/_2058_ ( .A(\mcsr/csr[2][13] ), .Z(\mcsr/_0196_ ) );
BUF_X1 \mcsr/_2059_ ( .A(\mcsr/_0806_ ), .Z(\csr_rdata[13] ) );
BUF_X1 \mcsr/_2060_ ( .A(\mcsr/csr[1][14] ), .Z(\mcsr/_0165_ ) );
BUF_X1 \mcsr/_2061_ ( .A(\mcsr/csr[0][14] ), .Z(\mcsr/_0133_ ) );
BUF_X1 \mcsr/_2062_ ( .A(\mcsr/csr[3][14] ), .Z(\mcsr/_0229_ ) );
BUF_X1 \mcsr/_2063_ ( .A(\mcsr/csr[2][14] ), .Z(\mcsr/_0197_ ) );
BUF_X1 \mcsr/_2064_ ( .A(\mcsr/_0807_ ), .Z(\csr_rdata[14] ) );
BUF_X1 \mcsr/_2065_ ( .A(\mcsr/csr[1][15] ), .Z(\mcsr/_0166_ ) );
BUF_X1 \mcsr/_2066_ ( .A(\mcsr/csr[0][15] ), .Z(\mcsr/_0134_ ) );
BUF_X1 \mcsr/_2067_ ( .A(\mcsr/csr[3][15] ), .Z(\mcsr/_0230_ ) );
BUF_X1 \mcsr/_2068_ ( .A(\mcsr/csr[2][15] ), .Z(\mcsr/_0198_ ) );
BUF_X1 \mcsr/_2069_ ( .A(\mcsr/_0808_ ), .Z(\csr_rdata[15] ) );
BUF_X1 \mcsr/_2070_ ( .A(\mcsr/csr[1][16] ), .Z(\mcsr/_0167_ ) );
BUF_X1 \mcsr/_2071_ ( .A(\mcsr/csr[0][16] ), .Z(\mcsr/_0135_ ) );
BUF_X1 \mcsr/_2072_ ( .A(\mcsr/csr[3][16] ), .Z(\mcsr/_0231_ ) );
BUF_X1 \mcsr/_2073_ ( .A(\mcsr/csr[2][16] ), .Z(\mcsr/_0199_ ) );
BUF_X1 \mcsr/_2074_ ( .A(\mcsr/_0809_ ), .Z(\csr_rdata[16] ) );
BUF_X1 \mcsr/_2075_ ( .A(\mcsr/csr[1][17] ), .Z(\mcsr/_0168_ ) );
BUF_X1 \mcsr/_2076_ ( .A(\mcsr/csr[0][17] ), .Z(\mcsr/_0136_ ) );
BUF_X1 \mcsr/_2077_ ( .A(\mcsr/csr[3][17] ), .Z(\mcsr/_0232_ ) );
BUF_X1 \mcsr/_2078_ ( .A(\mcsr/csr[2][17] ), .Z(\mcsr/_0200_ ) );
BUF_X1 \mcsr/_2079_ ( .A(\mcsr/_0810_ ), .Z(\csr_rdata[17] ) );
BUF_X1 \mcsr/_2080_ ( .A(\mcsr/csr[1][18] ), .Z(\mcsr/_0169_ ) );
BUF_X1 \mcsr/_2081_ ( .A(\mcsr/csr[0][18] ), .Z(\mcsr/_0137_ ) );
BUF_X1 \mcsr/_2082_ ( .A(\mcsr/csr[3][18] ), .Z(\mcsr/_0233_ ) );
BUF_X1 \mcsr/_2083_ ( .A(\mcsr/csr[2][18] ), .Z(\mcsr/_0201_ ) );
BUF_X1 \mcsr/_2084_ ( .A(\mcsr/_0811_ ), .Z(\csr_rdata[18] ) );
BUF_X1 \mcsr/_2085_ ( .A(\mcsr/csr[1][19] ), .Z(\mcsr/_0170_ ) );
BUF_X1 \mcsr/_2086_ ( .A(\mcsr/csr[0][19] ), .Z(\mcsr/_0138_ ) );
BUF_X1 \mcsr/_2087_ ( .A(\mcsr/csr[3][19] ), .Z(\mcsr/_0234_ ) );
BUF_X1 \mcsr/_2088_ ( .A(\mcsr/csr[2][19] ), .Z(\mcsr/_0202_ ) );
BUF_X1 \mcsr/_2089_ ( .A(\mcsr/_0812_ ), .Z(\csr_rdata[19] ) );
BUF_X1 \mcsr/_2090_ ( .A(\mcsr/csr[1][20] ), .Z(\mcsr/_0172_ ) );
BUF_X1 \mcsr/_2091_ ( .A(\mcsr/csr[0][20] ), .Z(\mcsr/_0140_ ) );
BUF_X1 \mcsr/_2092_ ( .A(\mcsr/csr[3][20] ), .Z(\mcsr/_0236_ ) );
BUF_X1 \mcsr/_2093_ ( .A(\mcsr/csr[2][20] ), .Z(\mcsr/_0204_ ) );
BUF_X1 \mcsr/_2094_ ( .A(\mcsr/_0814_ ), .Z(\csr_rdata[20] ) );
BUF_X1 \mcsr/_2095_ ( .A(\mcsr/csr[1][21] ), .Z(\mcsr/_0173_ ) );
BUF_X1 \mcsr/_2096_ ( .A(\mcsr/csr[0][21] ), .Z(\mcsr/_0141_ ) );
BUF_X1 \mcsr/_2097_ ( .A(\mcsr/csr[3][21] ), .Z(\mcsr/_0237_ ) );
BUF_X1 \mcsr/_2098_ ( .A(\mcsr/csr[2][21] ), .Z(\mcsr/_0205_ ) );
BUF_X1 \mcsr/_2099_ ( .A(\mcsr/_0815_ ), .Z(\csr_rdata[21] ) );
BUF_X1 \mcsr/_2100_ ( .A(\mcsr/csr[1][22] ), .Z(\mcsr/_0174_ ) );
BUF_X1 \mcsr/_2101_ ( .A(\mcsr/csr[0][22] ), .Z(\mcsr/_0142_ ) );
BUF_X1 \mcsr/_2102_ ( .A(\mcsr/csr[3][22] ), .Z(\mcsr/_0238_ ) );
BUF_X1 \mcsr/_2103_ ( .A(\mcsr/csr[2][22] ), .Z(\mcsr/_0206_ ) );
BUF_X1 \mcsr/_2104_ ( .A(\mcsr/_0816_ ), .Z(\csr_rdata[22] ) );
BUF_X1 \mcsr/_2105_ ( .A(\mcsr/csr[1][23] ), .Z(\mcsr/_0175_ ) );
BUF_X1 \mcsr/_2106_ ( .A(\mcsr/csr[0][23] ), .Z(\mcsr/_0143_ ) );
BUF_X1 \mcsr/_2107_ ( .A(\mcsr/csr[3][23] ), .Z(\mcsr/_0239_ ) );
BUF_X1 \mcsr/_2108_ ( .A(\mcsr/csr[2][23] ), .Z(\mcsr/_0207_ ) );
BUF_X1 \mcsr/_2109_ ( .A(\mcsr/_0817_ ), .Z(\csr_rdata[23] ) );
BUF_X1 \mcsr/_2110_ ( .A(\mcsr/csr[1][24] ), .Z(\mcsr/_0176_ ) );
BUF_X1 \mcsr/_2111_ ( .A(\mcsr/csr[0][24] ), .Z(\mcsr/_0144_ ) );
BUF_X1 \mcsr/_2112_ ( .A(\mcsr/csr[3][24] ), .Z(\mcsr/_0240_ ) );
BUF_X1 \mcsr/_2113_ ( .A(\mcsr/csr[2][24] ), .Z(\mcsr/_0208_ ) );
BUF_X1 \mcsr/_2114_ ( .A(\mcsr/_0818_ ), .Z(\csr_rdata[24] ) );
BUF_X1 \mcsr/_2115_ ( .A(\mcsr/csr[1][25] ), .Z(\mcsr/_0177_ ) );
BUF_X1 \mcsr/_2116_ ( .A(\mcsr/csr[0][25] ), .Z(\mcsr/_0145_ ) );
BUF_X1 \mcsr/_2117_ ( .A(\mcsr/csr[3][25] ), .Z(\mcsr/_0241_ ) );
BUF_X1 \mcsr/_2118_ ( .A(\mcsr/csr[2][25] ), .Z(\mcsr/_0209_ ) );
BUF_X1 \mcsr/_2119_ ( .A(\mcsr/_0819_ ), .Z(\csr_rdata[25] ) );
BUF_X1 \mcsr/_2120_ ( .A(\mcsr/csr[1][26] ), .Z(\mcsr/_0178_ ) );
BUF_X1 \mcsr/_2121_ ( .A(\mcsr/csr[0][26] ), .Z(\mcsr/_0146_ ) );
BUF_X1 \mcsr/_2122_ ( .A(\mcsr/csr[3][26] ), .Z(\mcsr/_0242_ ) );
BUF_X1 \mcsr/_2123_ ( .A(\mcsr/csr[2][26] ), .Z(\mcsr/_0210_ ) );
BUF_X1 \mcsr/_2124_ ( .A(\mcsr/_0820_ ), .Z(\csr_rdata[26] ) );
BUF_X1 \mcsr/_2125_ ( .A(\mcsr/csr[1][27] ), .Z(\mcsr/_0179_ ) );
BUF_X1 \mcsr/_2126_ ( .A(\mcsr/csr[0][27] ), .Z(\mcsr/_0147_ ) );
BUF_X1 \mcsr/_2127_ ( .A(\mcsr/csr[3][27] ), .Z(\mcsr/_0243_ ) );
BUF_X1 \mcsr/_2128_ ( .A(\mcsr/csr[2][27] ), .Z(\mcsr/_0211_ ) );
BUF_X1 \mcsr/_2129_ ( .A(\mcsr/_0821_ ), .Z(\csr_rdata[27] ) );
BUF_X1 \mcsr/_2130_ ( .A(\mcsr/csr[1][28] ), .Z(\mcsr/_0180_ ) );
BUF_X1 \mcsr/_2131_ ( .A(\mcsr/csr[0][28] ), .Z(\mcsr/_0148_ ) );
BUF_X1 \mcsr/_2132_ ( .A(\mcsr/csr[3][28] ), .Z(\mcsr/_0244_ ) );
BUF_X1 \mcsr/_2133_ ( .A(\mcsr/csr[2][28] ), .Z(\mcsr/_0212_ ) );
BUF_X1 \mcsr/_2134_ ( .A(\mcsr/_0822_ ), .Z(\csr_rdata[28] ) );
BUF_X1 \mcsr/_2135_ ( .A(\mcsr/csr[1][29] ), .Z(\mcsr/_0181_ ) );
BUF_X1 \mcsr/_2136_ ( .A(\mcsr/csr[0][29] ), .Z(\mcsr/_0149_ ) );
BUF_X1 \mcsr/_2137_ ( .A(\mcsr/csr[3][29] ), .Z(\mcsr/_0245_ ) );
BUF_X1 \mcsr/_2138_ ( .A(\mcsr/csr[2][29] ), .Z(\mcsr/_0213_ ) );
BUF_X1 \mcsr/_2139_ ( .A(\mcsr/_0823_ ), .Z(\csr_rdata[29] ) );
BUF_X1 \mcsr/_2140_ ( .A(\mcsr/csr[1][30] ), .Z(\mcsr/_0183_ ) );
BUF_X1 \mcsr/_2141_ ( .A(\mcsr/csr[0][30] ), .Z(\mcsr/_0151_ ) );
BUF_X1 \mcsr/_2142_ ( .A(\mcsr/csr[3][30] ), .Z(\mcsr/_0247_ ) );
BUF_X1 \mcsr/_2143_ ( .A(\mcsr/csr[2][30] ), .Z(\mcsr/_0215_ ) );
BUF_X1 \mcsr/_2144_ ( .A(\mcsr/_0825_ ), .Z(\csr_rdata[30] ) );
BUF_X1 \mcsr/_2145_ ( .A(\mcsr/csr[1][31] ), .Z(\mcsr/_0184_ ) );
BUF_X1 \mcsr/_2146_ ( .A(\mcsr/csr[0][31] ), .Z(\mcsr/_0152_ ) );
BUF_X1 \mcsr/_2147_ ( .A(\mcsr/csr[3][31] ), .Z(\mcsr/_0248_ ) );
BUF_X1 \mcsr/_2148_ ( .A(\mcsr/csr[2][31] ), .Z(\mcsr/_0216_ ) );
BUF_X1 \mcsr/_2149_ ( .A(\mcsr/_0826_ ), .Z(\csr_rdata[31] ) );
BUF_X1 \mcsr/_2150_ ( .A(\alu_result[0] ), .Z(\mcsr/_0866_ ) );
BUF_X1 \mcsr/_2151_ ( .A(\pc[0] ), .Z(\mcsr/_0770_ ) );
BUF_X1 \mcsr/_2152_ ( .A(\alu_result[1] ), .Z(\mcsr/_0877_ ) );
BUF_X1 \mcsr/_2153_ ( .A(\pc[1] ), .Z(\mcsr/_0781_ ) );
BUF_X1 \mcsr/_2154_ ( .A(\alu_result[2] ), .Z(\mcsr/_0888_ ) );
BUF_X1 \mcsr/_2155_ ( .A(\pc[2] ), .Z(\mcsr/_0792_ ) );
BUF_X1 \mcsr/_2156_ ( .A(\alu_result[3] ), .Z(\mcsr/_0891_ ) );
BUF_X1 \mcsr/_2157_ ( .A(\pc[3] ), .Z(\mcsr/_0795_ ) );
BUF_X1 \mcsr/_2158_ ( .A(\alu_result[4] ), .Z(\mcsr/_0892_ ) );
BUF_X1 \mcsr/_2159_ ( .A(\pc[4] ), .Z(\mcsr/_0796_ ) );
BUF_X1 \mcsr/_2160_ ( .A(\alu_result[5] ), .Z(\mcsr/_0893_ ) );
BUF_X1 \mcsr/_2161_ ( .A(\pc[5] ), .Z(\mcsr/_0797_ ) );
BUF_X1 \mcsr/_2162_ ( .A(\alu_result[6] ), .Z(\mcsr/_0894_ ) );
BUF_X1 \mcsr/_2163_ ( .A(\pc[6] ), .Z(\mcsr/_0798_ ) );
BUF_X1 \mcsr/_2164_ ( .A(\alu_result[7] ), .Z(\mcsr/_0895_ ) );
BUF_X1 \mcsr/_2165_ ( .A(\pc[7] ), .Z(\mcsr/_0799_ ) );
BUF_X1 \mcsr/_2166_ ( .A(\alu_result[8] ), .Z(\mcsr/_0896_ ) );
BUF_X1 \mcsr/_2167_ ( .A(\pc[8] ), .Z(\mcsr/_0800_ ) );
BUF_X1 \mcsr/_2168_ ( .A(\alu_result[9] ), .Z(\mcsr/_0897_ ) );
BUF_X1 \mcsr/_2169_ ( .A(\pc[9] ), .Z(\mcsr/_0801_ ) );
BUF_X1 \mcsr/_2170_ ( .A(\alu_result[10] ), .Z(\mcsr/_0867_ ) );
BUF_X1 \mcsr/_2171_ ( .A(\pc[10] ), .Z(\mcsr/_0771_ ) );
BUF_X1 \mcsr/_2172_ ( .A(\alu_result[11] ), .Z(\mcsr/_0868_ ) );
BUF_X1 \mcsr/_2173_ ( .A(\pc[11] ), .Z(\mcsr/_0772_ ) );
BUF_X1 \mcsr/_2174_ ( .A(\alu_result[12] ), .Z(\mcsr/_0869_ ) );
BUF_X1 \mcsr/_2175_ ( .A(\pc[12] ), .Z(\mcsr/_0773_ ) );
BUF_X1 \mcsr/_2176_ ( .A(\alu_result[13] ), .Z(\mcsr/_0870_ ) );
BUF_X1 \mcsr/_2177_ ( .A(\pc[13] ), .Z(\mcsr/_0774_ ) );
BUF_X1 \mcsr/_2178_ ( .A(\alu_result[14] ), .Z(\mcsr/_0871_ ) );
BUF_X1 \mcsr/_2179_ ( .A(\pc[14] ), .Z(\mcsr/_0775_ ) );
BUF_X1 \mcsr/_2180_ ( .A(\alu_result[15] ), .Z(\mcsr/_0872_ ) );
BUF_X1 \mcsr/_2181_ ( .A(\pc[15] ), .Z(\mcsr/_0776_ ) );
BUF_X1 \mcsr/_2182_ ( .A(\alu_result[16] ), .Z(\mcsr/_0873_ ) );
BUF_X1 \mcsr/_2183_ ( .A(\pc[16] ), .Z(\mcsr/_0777_ ) );
BUF_X1 \mcsr/_2184_ ( .A(\alu_result[17] ), .Z(\mcsr/_0874_ ) );
BUF_X1 \mcsr/_2185_ ( .A(\pc[17] ), .Z(\mcsr/_0778_ ) );
BUF_X1 \mcsr/_2186_ ( .A(\alu_result[18] ), .Z(\mcsr/_0875_ ) );
BUF_X1 \mcsr/_2187_ ( .A(\pc[18] ), .Z(\mcsr/_0779_ ) );
BUF_X1 \mcsr/_2188_ ( .A(\alu_result[19] ), .Z(\mcsr/_0876_ ) );
BUF_X1 \mcsr/_2189_ ( .A(\pc[19] ), .Z(\mcsr/_0780_ ) );
BUF_X1 \mcsr/_2190_ ( .A(\alu_result[20] ), .Z(\mcsr/_0878_ ) );
BUF_X1 \mcsr/_2191_ ( .A(\pc[20] ), .Z(\mcsr/_0782_ ) );
BUF_X1 \mcsr/_2192_ ( .A(\alu_result[21] ), .Z(\mcsr/_0879_ ) );
BUF_X1 \mcsr/_2193_ ( .A(\pc[21] ), .Z(\mcsr/_0783_ ) );
BUF_X1 \mcsr/_2194_ ( .A(\alu_result[22] ), .Z(\mcsr/_0880_ ) );
BUF_X1 \mcsr/_2195_ ( .A(\pc[22] ), .Z(\mcsr/_0784_ ) );
BUF_X1 \mcsr/_2196_ ( .A(\alu_result[23] ), .Z(\mcsr/_0881_ ) );
BUF_X1 \mcsr/_2197_ ( .A(\pc[23] ), .Z(\mcsr/_0785_ ) );
BUF_X1 \mcsr/_2198_ ( .A(\alu_result[24] ), .Z(\mcsr/_0882_ ) );
BUF_X1 \mcsr/_2199_ ( .A(\pc[24] ), .Z(\mcsr/_0786_ ) );
BUF_X1 \mcsr/_2200_ ( .A(\alu_result[25] ), .Z(\mcsr/_0883_ ) );
BUF_X1 \mcsr/_2201_ ( .A(\pc[25] ), .Z(\mcsr/_0787_ ) );
BUF_X1 \mcsr/_2202_ ( .A(\alu_result[26] ), .Z(\mcsr/_0884_ ) );
BUF_X1 \mcsr/_2203_ ( .A(\pc[26] ), .Z(\mcsr/_0788_ ) );
BUF_X1 \mcsr/_2204_ ( .A(\alu_result[27] ), .Z(\mcsr/_0885_ ) );
BUF_X1 \mcsr/_2205_ ( .A(\pc[27] ), .Z(\mcsr/_0789_ ) );
BUF_X1 \mcsr/_2206_ ( .A(\alu_result[28] ), .Z(\mcsr/_0886_ ) );
BUF_X1 \mcsr/_2207_ ( .A(\pc[28] ), .Z(\mcsr/_0790_ ) );
BUF_X1 \mcsr/_2208_ ( .A(\alu_result[29] ), .Z(\mcsr/_0887_ ) );
BUF_X1 \mcsr/_2209_ ( .A(\pc[29] ), .Z(\mcsr/_0791_ ) );
BUF_X1 \mcsr/_2210_ ( .A(\alu_result[30] ), .Z(\mcsr/_0889_ ) );
BUF_X1 \mcsr/_2211_ ( .A(\pc[30] ), .Z(\mcsr/_0793_ ) );
BUF_X1 \mcsr/_2212_ ( .A(\alu_result[31] ), .Z(\mcsr/_0890_ ) );
BUF_X1 \mcsr/_2213_ ( .A(\pc[31] ), .Z(\mcsr/_0794_ ) );
BUF_X1 \mcsr/_2214_ ( .A(\mcsr/_0834_ ), .Z(\csr_upc[0] ) );
BUF_X1 \mcsr/_2215_ ( .A(\mcsr/_0845_ ), .Z(\csr_upc[1] ) );
BUF_X1 \mcsr/_2216_ ( .A(\mcsr/_0856_ ), .Z(\csr_upc[2] ) );
BUF_X1 \mcsr/_2217_ ( .A(\mcsr/_0859_ ), .Z(\csr_upc[3] ) );
BUF_X1 \mcsr/_2218_ ( .A(\mcsr/_0860_ ), .Z(\csr_upc[4] ) );
BUF_X1 \mcsr/_2219_ ( .A(\mcsr/_0861_ ), .Z(\csr_upc[5] ) );
BUF_X1 \mcsr/_2220_ ( .A(\mcsr/_0862_ ), .Z(\csr_upc[6] ) );
BUF_X1 \mcsr/_2221_ ( .A(\mcsr/_0863_ ), .Z(\csr_upc[7] ) );
BUF_X1 \mcsr/_2222_ ( .A(\mcsr/_0864_ ), .Z(\csr_upc[8] ) );
BUF_X1 \mcsr/_2223_ ( .A(\mcsr/_0865_ ), .Z(\csr_upc[9] ) );
BUF_X1 \mcsr/_2224_ ( .A(\mcsr/_0835_ ), .Z(\csr_upc[10] ) );
BUF_X1 \mcsr/_2225_ ( .A(\mcsr/_0836_ ), .Z(\csr_upc[11] ) );
BUF_X1 \mcsr/_2226_ ( .A(\mcsr/_0837_ ), .Z(\csr_upc[12] ) );
BUF_X1 \mcsr/_2227_ ( .A(\mcsr/_0838_ ), .Z(\csr_upc[13] ) );
BUF_X1 \mcsr/_2228_ ( .A(\mcsr/_0839_ ), .Z(\csr_upc[14] ) );
BUF_X1 \mcsr/_2229_ ( .A(\mcsr/_0840_ ), .Z(\csr_upc[15] ) );
BUF_X1 \mcsr/_2230_ ( .A(\mcsr/_0841_ ), .Z(\csr_upc[16] ) );
BUF_X1 \mcsr/_2231_ ( .A(\mcsr/_0842_ ), .Z(\csr_upc[17] ) );
BUF_X1 \mcsr/_2232_ ( .A(\mcsr/_0843_ ), .Z(\csr_upc[18] ) );
BUF_X1 \mcsr/_2233_ ( .A(\mcsr/_0844_ ), .Z(\csr_upc[19] ) );
BUF_X1 \mcsr/_2234_ ( .A(\mcsr/_0846_ ), .Z(\csr_upc[20] ) );
BUF_X1 \mcsr/_2235_ ( .A(\mcsr/_0847_ ), .Z(\csr_upc[21] ) );
BUF_X1 \mcsr/_2236_ ( .A(\mcsr/_0848_ ), .Z(\csr_upc[22] ) );
BUF_X1 \mcsr/_2237_ ( .A(\mcsr/_0849_ ), .Z(\csr_upc[23] ) );
BUF_X1 \mcsr/_2238_ ( .A(\mcsr/_0850_ ), .Z(\csr_upc[24] ) );
BUF_X1 \mcsr/_2239_ ( .A(\mcsr/_0851_ ), .Z(\csr_upc[25] ) );
BUF_X1 \mcsr/_2240_ ( .A(\mcsr/_0852_ ), .Z(\csr_upc[26] ) );
BUF_X1 \mcsr/_2241_ ( .A(\mcsr/_0853_ ), .Z(\csr_upc[27] ) );
BUF_X1 \mcsr/_2242_ ( .A(\mcsr/_0854_ ), .Z(\csr_upc[28] ) );
BUF_X1 \mcsr/_2243_ ( .A(\mcsr/_0855_ ), .Z(\csr_upc[29] ) );
BUF_X1 \mcsr/_2244_ ( .A(\mcsr/_0857_ ), .Z(\csr_upc[30] ) );
BUF_X1 \mcsr/_2245_ ( .A(\mcsr/_0858_ ), .Z(\csr_upc[31] ) );
BUF_X1 \mcsr/_2246_ ( .A(\mcsr/_0000_ ), .Z(\mcsr/_1027_ ) );
BUF_X1 \mcsr/_2247_ ( .A(\mcsr/_0001_ ), .Z(\mcsr/_1028_ ) );
BUF_X1 \mcsr/_2248_ ( .A(\mcsr/_0002_ ), .Z(\mcsr/_1029_ ) );
BUF_X1 \mcsr/_2249_ ( .A(\mcsr/_0003_ ), .Z(\mcsr/_1030_ ) );
BUF_X1 \mcsr/_2250_ ( .A(\mcsr/_0004_ ), .Z(\mcsr/_1031_ ) );
BUF_X1 \mcsr/_2251_ ( .A(\mcsr/_0005_ ), .Z(\mcsr/_1032_ ) );
BUF_X1 \mcsr/_2252_ ( .A(\mcsr/_0006_ ), .Z(\mcsr/_1033_ ) );
BUF_X1 \mcsr/_2253_ ( .A(\mcsr/_0007_ ), .Z(\mcsr/_1034_ ) );
BUF_X1 \mcsr/_2254_ ( .A(\mcsr/_0008_ ), .Z(\mcsr/_1035_ ) );
BUF_X1 \mcsr/_2255_ ( .A(\mcsr/_0009_ ), .Z(\mcsr/_1036_ ) );
BUF_X1 \mcsr/_2256_ ( .A(\mcsr/_0010_ ), .Z(\mcsr/_1037_ ) );
BUF_X1 \mcsr/_2257_ ( .A(\mcsr/_0011_ ), .Z(\mcsr/_1038_ ) );
BUF_X1 \mcsr/_2258_ ( .A(\mcsr/_0012_ ), .Z(\mcsr/_1039_ ) );
BUF_X1 \mcsr/_2259_ ( .A(\mcsr/_0013_ ), .Z(\mcsr/_1040_ ) );
BUF_X1 \mcsr/_2260_ ( .A(\mcsr/_0014_ ), .Z(\mcsr/_1041_ ) );
BUF_X1 \mcsr/_2261_ ( .A(\mcsr/_0015_ ), .Z(\mcsr/_1042_ ) );
BUF_X1 \mcsr/_2262_ ( .A(\mcsr/_0016_ ), .Z(\mcsr/_1043_ ) );
BUF_X1 \mcsr/_2263_ ( .A(\mcsr/_0017_ ), .Z(\mcsr/_1044_ ) );
BUF_X1 \mcsr/_2264_ ( .A(\mcsr/_0018_ ), .Z(\mcsr/_1045_ ) );
BUF_X1 \mcsr/_2265_ ( .A(\mcsr/_0019_ ), .Z(\mcsr/_1046_ ) );
BUF_X1 \mcsr/_2266_ ( .A(\mcsr/_0020_ ), .Z(\mcsr/_1047_ ) );
BUF_X1 \mcsr/_2267_ ( .A(\mcsr/_0021_ ), .Z(\mcsr/_1048_ ) );
BUF_X1 \mcsr/_2268_ ( .A(\mcsr/_0022_ ), .Z(\mcsr/_1049_ ) );
BUF_X1 \mcsr/_2269_ ( .A(\mcsr/_0023_ ), .Z(\mcsr/_1050_ ) );
BUF_X1 \mcsr/_2270_ ( .A(\mcsr/_0024_ ), .Z(\mcsr/_1051_ ) );
BUF_X1 \mcsr/_2271_ ( .A(\mcsr/_0025_ ), .Z(\mcsr/_1052_ ) );
BUF_X1 \mcsr/_2272_ ( .A(\mcsr/_0026_ ), .Z(\mcsr/_1053_ ) );
BUF_X1 \mcsr/_2273_ ( .A(\mcsr/_0027_ ), .Z(\mcsr/_1054_ ) );
BUF_X1 \mcsr/_2274_ ( .A(\mcsr/_0028_ ), .Z(\mcsr/_1055_ ) );
BUF_X1 \mcsr/_2275_ ( .A(\mcsr/_0029_ ), .Z(\mcsr/_1056_ ) );
BUF_X1 \mcsr/_2276_ ( .A(\mcsr/_0030_ ), .Z(\mcsr/_1057_ ) );
BUF_X1 \mcsr/_2277_ ( .A(\mcsr/_0031_ ), .Z(\mcsr/_1058_ ) );
BUF_X1 \mcsr/_2278_ ( .A(\mcsr/_0032_ ), .Z(\mcsr/_1059_ ) );
BUF_X1 \mcsr/_2279_ ( .A(\mcsr/_0033_ ), .Z(\mcsr/_1060_ ) );
BUF_X1 \mcsr/_2280_ ( .A(\mcsr/_0034_ ), .Z(\mcsr/_1061_ ) );
BUF_X1 \mcsr/_2281_ ( .A(\mcsr/_0035_ ), .Z(\mcsr/_1062_ ) );
BUF_X1 \mcsr/_2282_ ( .A(\mcsr/_0036_ ), .Z(\mcsr/_1063_ ) );
BUF_X1 \mcsr/_2283_ ( .A(\mcsr/_0037_ ), .Z(\mcsr/_1064_ ) );
BUF_X1 \mcsr/_2284_ ( .A(\mcsr/_0038_ ), .Z(\mcsr/_1065_ ) );
BUF_X1 \mcsr/_2285_ ( .A(\mcsr/_0039_ ), .Z(\mcsr/_1066_ ) );
BUF_X1 \mcsr/_2286_ ( .A(\mcsr/_0040_ ), .Z(\mcsr/_1067_ ) );
BUF_X1 \mcsr/_2287_ ( .A(\mcsr/_0041_ ), .Z(\mcsr/_1068_ ) );
BUF_X1 \mcsr/_2288_ ( .A(\mcsr/_0042_ ), .Z(\mcsr/_1069_ ) );
BUF_X1 \mcsr/_2289_ ( .A(\mcsr/_0043_ ), .Z(\mcsr/_1070_ ) );
BUF_X1 \mcsr/_2290_ ( .A(\mcsr/_0044_ ), .Z(\mcsr/_1071_ ) );
BUF_X1 \mcsr/_2291_ ( .A(\mcsr/_0045_ ), .Z(\mcsr/_1072_ ) );
BUF_X1 \mcsr/_2292_ ( .A(\mcsr/_0046_ ), .Z(\mcsr/_1073_ ) );
BUF_X1 \mcsr/_2293_ ( .A(\mcsr/_0047_ ), .Z(\mcsr/_1074_ ) );
BUF_X1 \mcsr/_2294_ ( .A(\mcsr/_0048_ ), .Z(\mcsr/_1075_ ) );
BUF_X1 \mcsr/_2295_ ( .A(\mcsr/_0049_ ), .Z(\mcsr/_1076_ ) );
BUF_X1 \mcsr/_2296_ ( .A(\mcsr/_0050_ ), .Z(\mcsr/_1077_ ) );
BUF_X1 \mcsr/_2297_ ( .A(\mcsr/_0051_ ), .Z(\mcsr/_1078_ ) );
BUF_X1 \mcsr/_2298_ ( .A(\mcsr/_0052_ ), .Z(\mcsr/_1079_ ) );
BUF_X1 \mcsr/_2299_ ( .A(\mcsr/_0053_ ), .Z(\mcsr/_1080_ ) );
BUF_X1 \mcsr/_2300_ ( .A(\mcsr/_0054_ ), .Z(\mcsr/_1081_ ) );
BUF_X1 \mcsr/_2301_ ( .A(\mcsr/_0055_ ), .Z(\mcsr/_1082_ ) );
BUF_X1 \mcsr/_2302_ ( .A(\mcsr/_0056_ ), .Z(\mcsr/_1083_ ) );
BUF_X1 \mcsr/_2303_ ( .A(\mcsr/_0057_ ), .Z(\mcsr/_1084_ ) );
BUF_X1 \mcsr/_2304_ ( .A(\mcsr/_0058_ ), .Z(\mcsr/_1085_ ) );
BUF_X1 \mcsr/_2305_ ( .A(\mcsr/_0059_ ), .Z(\mcsr/_1086_ ) );
BUF_X1 \mcsr/_2306_ ( .A(\mcsr/_0060_ ), .Z(\mcsr/_1087_ ) );
BUF_X1 \mcsr/_2307_ ( .A(\mcsr/_0061_ ), .Z(\mcsr/_1088_ ) );
BUF_X1 \mcsr/_2308_ ( .A(\mcsr/_0062_ ), .Z(\mcsr/_1089_ ) );
BUF_X1 \mcsr/_2309_ ( .A(\mcsr/_0063_ ), .Z(\mcsr/_1090_ ) );
BUF_X1 \mcsr/_2310_ ( .A(\mcsr/_0096_ ), .Z(\mcsr/_1123_ ) );
BUF_X1 \mcsr/_2311_ ( .A(\mcsr/_0097_ ), .Z(\mcsr/_1124_ ) );
BUF_X1 \mcsr/_2312_ ( .A(\mcsr/_0098_ ), .Z(\mcsr/_1125_ ) );
BUF_X1 \mcsr/_2313_ ( .A(\mcsr/_0099_ ), .Z(\mcsr/_1126_ ) );
BUF_X1 \mcsr/_2314_ ( .A(\mcsr/_0100_ ), .Z(\mcsr/_1127_ ) );
BUF_X1 \mcsr/_2315_ ( .A(\mcsr/_0101_ ), .Z(\mcsr/_1128_ ) );
BUF_X1 \mcsr/_2316_ ( .A(\mcsr/_0102_ ), .Z(\mcsr/_1129_ ) );
BUF_X1 \mcsr/_2317_ ( .A(\mcsr/_0103_ ), .Z(\mcsr/_1130_ ) );
BUF_X1 \mcsr/_2318_ ( .A(\mcsr/_0104_ ), .Z(\mcsr/_1131_ ) );
BUF_X1 \mcsr/_2319_ ( .A(\mcsr/_0105_ ), .Z(\mcsr/_1132_ ) );
BUF_X1 \mcsr/_2320_ ( .A(\mcsr/_0106_ ), .Z(\mcsr/_1133_ ) );
BUF_X1 \mcsr/_2321_ ( .A(\mcsr/_0107_ ), .Z(\mcsr/_1134_ ) );
BUF_X1 \mcsr/_2322_ ( .A(\mcsr/_0108_ ), .Z(\mcsr/_1135_ ) );
BUF_X1 \mcsr/_2323_ ( .A(\mcsr/_0109_ ), .Z(\mcsr/_1136_ ) );
BUF_X1 \mcsr/_2324_ ( .A(\mcsr/_0110_ ), .Z(\mcsr/_1137_ ) );
BUF_X1 \mcsr/_2325_ ( .A(\mcsr/_0111_ ), .Z(\mcsr/_1138_ ) );
BUF_X1 \mcsr/_2326_ ( .A(\mcsr/_0112_ ), .Z(\mcsr/_1139_ ) );
BUF_X1 \mcsr/_2327_ ( .A(\mcsr/_0113_ ), .Z(\mcsr/_1140_ ) );
BUF_X1 \mcsr/_2328_ ( .A(\mcsr/_0114_ ), .Z(\mcsr/_1141_ ) );
BUF_X1 \mcsr/_2329_ ( .A(\mcsr/_0115_ ), .Z(\mcsr/_1142_ ) );
BUF_X1 \mcsr/_2330_ ( .A(\mcsr/_0116_ ), .Z(\mcsr/_1143_ ) );
BUF_X1 \mcsr/_2331_ ( .A(\mcsr/_0117_ ), .Z(\mcsr/_1144_ ) );
BUF_X1 \mcsr/_2332_ ( .A(\mcsr/_0118_ ), .Z(\mcsr/_1145_ ) );
BUF_X1 \mcsr/_2333_ ( .A(\mcsr/_0119_ ), .Z(\mcsr/_1146_ ) );
BUF_X1 \mcsr/_2334_ ( .A(\mcsr/_0120_ ), .Z(\mcsr/_1147_ ) );
BUF_X1 \mcsr/_2335_ ( .A(\mcsr/_0121_ ), .Z(\mcsr/_1148_ ) );
BUF_X1 \mcsr/_2336_ ( .A(\mcsr/_0122_ ), .Z(\mcsr/_1149_ ) );
BUF_X1 \mcsr/_2337_ ( .A(\mcsr/_0123_ ), .Z(\mcsr/_1150_ ) );
BUF_X1 \mcsr/_2338_ ( .A(\mcsr/_0124_ ), .Z(\mcsr/_1151_ ) );
BUF_X1 \mcsr/_2339_ ( .A(\mcsr/_0125_ ), .Z(\mcsr/_1152_ ) );
BUF_X1 \mcsr/_2340_ ( .A(\mcsr/_0126_ ), .Z(\mcsr/_1153_ ) );
BUF_X1 \mcsr/_2341_ ( .A(\mcsr/_0127_ ), .Z(\mcsr/_1154_ ) );
BUF_X1 \mcsr/_2342_ ( .A(\mcsr/_0064_ ), .Z(\mcsr/_1091_ ) );
BUF_X1 \mcsr/_2343_ ( .A(\mcsr/_0065_ ), .Z(\mcsr/_1092_ ) );
BUF_X1 \mcsr/_2344_ ( .A(\mcsr/_0066_ ), .Z(\mcsr/_1093_ ) );
BUF_X1 \mcsr/_2345_ ( .A(\mcsr/_0067_ ), .Z(\mcsr/_1094_ ) );
BUF_X1 \mcsr/_2346_ ( .A(\mcsr/_0068_ ), .Z(\mcsr/_1095_ ) );
BUF_X1 \mcsr/_2347_ ( .A(\mcsr/_0069_ ), .Z(\mcsr/_1096_ ) );
BUF_X1 \mcsr/_2348_ ( .A(\mcsr/_0070_ ), .Z(\mcsr/_1097_ ) );
BUF_X1 \mcsr/_2349_ ( .A(\mcsr/_0071_ ), .Z(\mcsr/_1098_ ) );
BUF_X1 \mcsr/_2350_ ( .A(\mcsr/_0072_ ), .Z(\mcsr/_1099_ ) );
BUF_X1 \mcsr/_2351_ ( .A(\mcsr/_0073_ ), .Z(\mcsr/_1100_ ) );
BUF_X1 \mcsr/_2352_ ( .A(\mcsr/_0074_ ), .Z(\mcsr/_1101_ ) );
BUF_X1 \mcsr/_2353_ ( .A(\mcsr/_0075_ ), .Z(\mcsr/_1102_ ) );
BUF_X1 \mcsr/_2354_ ( .A(\mcsr/_0076_ ), .Z(\mcsr/_1103_ ) );
BUF_X1 \mcsr/_2355_ ( .A(\mcsr/_0077_ ), .Z(\mcsr/_1104_ ) );
BUF_X1 \mcsr/_2356_ ( .A(\mcsr/_0078_ ), .Z(\mcsr/_1105_ ) );
BUF_X1 \mcsr/_2357_ ( .A(\mcsr/_0079_ ), .Z(\mcsr/_1106_ ) );
BUF_X1 \mcsr/_2358_ ( .A(\mcsr/_0080_ ), .Z(\mcsr/_1107_ ) );
BUF_X1 \mcsr/_2359_ ( .A(\mcsr/_0081_ ), .Z(\mcsr/_1108_ ) );
BUF_X1 \mcsr/_2360_ ( .A(\mcsr/_0082_ ), .Z(\mcsr/_1109_ ) );
BUF_X1 \mcsr/_2361_ ( .A(\mcsr/_0083_ ), .Z(\mcsr/_1110_ ) );
BUF_X1 \mcsr/_2362_ ( .A(\mcsr/_0084_ ), .Z(\mcsr/_1111_ ) );
BUF_X1 \mcsr/_2363_ ( .A(\mcsr/_0085_ ), .Z(\mcsr/_1112_ ) );
BUF_X1 \mcsr/_2364_ ( .A(\mcsr/_0086_ ), .Z(\mcsr/_1113_ ) );
BUF_X1 \mcsr/_2365_ ( .A(\mcsr/_0087_ ), .Z(\mcsr/_1114_ ) );
BUF_X1 \mcsr/_2366_ ( .A(\mcsr/_0088_ ), .Z(\mcsr/_1115_ ) );
BUF_X1 \mcsr/_2367_ ( .A(\mcsr/_0089_ ), .Z(\mcsr/_1116_ ) );
BUF_X1 \mcsr/_2368_ ( .A(\mcsr/_0090_ ), .Z(\mcsr/_1117_ ) );
BUF_X1 \mcsr/_2369_ ( .A(\mcsr/_0091_ ), .Z(\mcsr/_1118_ ) );
BUF_X1 \mcsr/_2370_ ( .A(\mcsr/_0092_ ), .Z(\mcsr/_1119_ ) );
BUF_X1 \mcsr/_2371_ ( .A(\mcsr/_0093_ ), .Z(\mcsr/_1120_ ) );
BUF_X1 \mcsr/_2372_ ( .A(\mcsr/_0094_ ), .Z(\mcsr/_1121_ ) );
BUF_X1 \mcsr/_2373_ ( .A(\mcsr/_0095_ ), .Z(\mcsr/_1122_ ) );
INV_X1 \mexu/_1094_ ( .A(\mexu/_0974_ ), .ZN(\mexu/_0365_ ) );
AND3_X1 \mexu/_1095_ ( .A1(\mexu/_0365_ ), .A2(\mexu/_0972_ ), .A3(\mexu/_0971_ ), .ZN(\mexu/_0366_ ) );
INV_X1 \mexu/_1096_ ( .A(\mexu/_0973_ ), .ZN(\mexu/_0367_ ) );
AND2_X2 \mexu/_1097_ ( .A1(\mexu/_0366_ ), .A2(\mexu/_0367_ ), .ZN(\mexu/_0368_ ) );
INV_X1 \mexu/_1098_ ( .A(\mexu/_0368_ ), .ZN(\mexu/_0369_ ) );
OR3_X1 \mexu/_1099_ ( .A1(\mexu/_0975_ ), .A2(\mexu/_0976_ ), .A3(\mexu/_0977_ ), .ZN(\mexu/_0370_ ) );
NOR2_X1 \mexu/_1100_ ( .A1(\mexu/_0369_ ), .A2(\mexu/_0370_ ), .ZN(\mexu/_0212_ ) );
AND3_X1 \mexu/_1101_ ( .A1(\mexu/_0975_ ), .A2(\mexu/_0976_ ), .A3(\mexu/_0977_ ), .ZN(\mexu/_0371_ ) );
BUF_X4 \mexu/_1102_ ( .A(\mexu/_0371_ ), .Z(\mexu/_0372_ ) );
AND2_X1 \mexu/_1103_ ( .A1(\mexu/_0368_ ), .A2(\mexu/_0372_ ), .ZN(\mexu/_0075_ ) );
BUF_X2 \mexu/_1104_ ( .A(\mexu/_0368_ ), .Z(\mexu/_0373_ ) );
BUF_X2 \mexu/_1105_ ( .A(\mexu/_0372_ ), .Z(\mexu/_0374_ ) );
NOR2_X1 \mexu/_1106_ ( .A1(\mexu/_0173_ ), .A2(\mexu/_0174_ ), .ZN(\mexu/_0375_ ) );
INV_X1 \mexu/_1107_ ( .A(\mexu/_0175_ ), .ZN(\mexu/_0376_ ) );
AND2_X2 \mexu/_1108_ ( .A1(\mexu/_0375_ ), .A2(\mexu/_0376_ ), .ZN(\mexu/_0377_ ) );
BUF_X2 \mexu/_1109_ ( .A(\mexu/_0377_ ), .Z(\mexu/_0378_ ) );
AND3_X1 \mexu/_1110_ ( .A1(\mexu/_0373_ ), .A2(\mexu/_0374_ ), .A3(\mexu/_0378_ ), .ZN(\mexu/_1085_ ) );
INV_X1 \mexu/_1111_ ( .A(\mexu/_0212_ ), .ZN(\mexu/_0379_ ) );
AND2_X1 \mexu/_1112_ ( .A1(\mexu/_0972_ ), .A2(\mexu/_0971_ ), .ZN(\mexu/_0380_ ) );
AND3_X1 \mexu/_1113_ ( .A1(\mexu/_0380_ ), .A2(\mexu/_0973_ ), .A3(\mexu/_0365_ ), .ZN(\mexu/_0381_ ) );
INV_X1 \mexu/_1114_ ( .A(\mexu/_0977_ ), .ZN(\mexu/_0382_ ) );
AND3_X1 \mexu/_1115_ ( .A1(\mexu/_0382_ ), .A2(\mexu/_0975_ ), .A3(\mexu/_0976_ ), .ZN(\mexu/_0383_ ) );
NAND2_X2 \mexu/_1116_ ( .A1(\mexu/_0381_ ), .A2(\mexu/_0383_ ), .ZN(\mexu/_0384_ ) );
AND2_X1 \mexu/_1117_ ( .A1(\mexu/_0379_ ), .A2(\mexu/_0384_ ), .ZN(\mexu/_0385_ ) );
INV_X1 \mexu/_1118_ ( .A(\mexu/_0975_ ), .ZN(\mexu/_0386_ ) );
AND3_X2 \mexu/_1119_ ( .A1(\mexu/_0386_ ), .A2(\mexu/_0976_ ), .A3(\mexu/_0977_ ), .ZN(\mexu/_0387_ ) );
AND2_X1 \mexu/_1120_ ( .A1(\mexu/_0381_ ), .A2(\mexu/_0387_ ), .ZN(\mexu/_0388_ ) );
AND4_X1 \mexu/_1121_ ( .A1(\mexu/_0972_ ), .A2(\mexu/_0971_ ), .A3(\mexu/_0973_ ), .A4(\mexu/_0974_ ), .ZN(\mexu/_0389_ ) );
AND2_X1 \mexu/_1122_ ( .A1(\mexu/_0387_ ), .A2(\mexu/_0389_ ), .ZN(\mexu/_0390_ ) );
NOR2_X2 \mexu/_1123_ ( .A1(\mexu/_0388_ ), .A2(\mexu/_0390_ ), .ZN(\mexu/_0391_ ) );
NOR3_X1 \mexu/_1124_ ( .A1(\mexu/_0386_ ), .A2(\mexu/_0976_ ), .A3(\mexu/_0977_ ), .ZN(\mexu/_0392_ ) );
AND2_X1 \mexu/_1125_ ( .A1(\mexu/_0381_ ), .A2(\mexu/_0392_ ), .ZN(\mexu/_0393_ ) );
BUF_X4 \mexu/_1126_ ( .A(\mexu/_0393_ ), .Z(\mexu/_0394_ ) );
INV_X2 \mexu/_1127_ ( .A(\mexu/_0394_ ), .ZN(\mexu/_0395_ ) );
AND2_X1 \mexu/_1128_ ( .A1(\mexu/_0391_ ), .A2(\mexu/_0395_ ), .ZN(\mexu/_0396_ ) );
INV_X1 \mexu/_1129_ ( .A(\mexu/_0075_ ), .ZN(\mexu/_0397_ ) );
AND2_X1 \mexu/_1130_ ( .A1(\mexu/_0366_ ), .A2(\mexu/_0392_ ), .ZN(\mexu/_0398_ ) );
AND2_X2 \mexu/_1131_ ( .A1(\mexu/_0398_ ), .A2(\mexu/_0367_ ), .ZN(\mexu/_0399_ ) );
AND2_X1 \mexu/_1132_ ( .A1(\mexu/_0368_ ), .A2(\mexu/_0383_ ), .ZN(\mexu/_0400_ ) );
NOR2_X1 \mexu/_1133_ ( .A1(\mexu/_0399_ ), .A2(\mexu/_0400_ ), .ZN(\mexu/_0401_ ) );
NAND4_X1 \mexu/_1134_ ( .A1(\mexu/_0385_ ), .A2(\mexu/_0396_ ), .A3(\mexu/_0397_ ), .A4(\mexu/_0401_ ), .ZN(\mexu/_1017_ ) );
NAND3_X1 \mexu/_1135_ ( .A1(\mexu/_0386_ ), .A2(\mexu/_0382_ ), .A3(\mexu/_0976_ ), .ZN(\mexu/_0402_ ) );
NOR2_X1 \mexu/_1136_ ( .A1(\mexu/_0369_ ), .A2(\mexu/_0402_ ), .ZN(\mexu/_0213_ ) );
AND2_X1 \mexu/_1137_ ( .A1(\mexu/_0368_ ), .A2(\mexu/_0387_ ), .ZN(\mexu/_0403_ ) );
OR2_X1 \mexu/_1138_ ( .A1(\mexu/_1017_ ), .A2(\mexu/_0403_ ), .ZN(\mexu/_0073_ ) );
INV_X1 \mexu/_1139_ ( .A(\mexu/_0173_ ), .ZN(\mexu/_0404_ ) );
NOR2_X1 \mexu/_1140_ ( .A1(\mexu/_0404_ ), .A2(\mexu/_0174_ ), .ZN(\mexu/_0405_ ) );
INV_X1 \mexu/_1141_ ( .A(\mexu/_0174_ ), .ZN(\mexu/_0406_ ) );
OAI21_X1 \mexu/_1142_ ( .A(\mexu/_0175_ ), .B1(\mexu/_0406_ ), .B2(\mexu/_0173_ ), .ZN(\mexu/_0407_ ) );
OR3_X1 \mexu/_1143_ ( .A1(\mexu/_0401_ ), .A2(\mexu/_0405_ ), .A3(\mexu/_0407_ ), .ZN(\mexu/_0408_ ) );
NOR2_X1 \mexu/_1144_ ( .A1(\mexu/_0406_ ), .A2(\mexu/_0175_ ), .ZN(\mexu/_0409_ ) );
INV_X1 \mexu/_1145_ ( .A(\mexu/_0409_ ), .ZN(\mexu/_0410_ ) );
AND3_X1 \mexu/_1146_ ( .A1(\mexu/_0368_ ), .A2(\mexu/_0387_ ), .A3(\mexu/_0410_ ), .ZN(\mexu/_0411_ ) );
INV_X1 \mexu/_1147_ ( .A(\mexu/_0411_ ), .ZN(\mexu/_0412_ ) );
AND2_X1 \mexu/_1148_ ( .A1(\mexu/_0405_ ), .A2(\mexu/_0175_ ), .ZN(\mexu/_0413_ ) );
INV_X1 \mexu/_1149_ ( .A(\mexu/_0413_ ), .ZN(\mexu/_0414_ ) );
INV_X1 \mexu/_1150_ ( .A(\mexu/_0203_ ), .ZN(\mexu/_0415_ ) );
BUF_X4 \mexu/_1151_ ( .A(\mexu/_0399_ ), .Z(\mexu/_0416_ ) );
INV_X1 \mexu/_1152_ ( .A(\mexu/_0177_ ), .ZN(\mexu/_0417_ ) );
AOI22_X1 \mexu/_1153_ ( .A1(\mexu/_0415_ ), .A2(\mexu/_0400_ ), .B1(\mexu/_0416_ ), .B2(\mexu/_0417_ ), .ZN(\mexu/_0418_ ) );
OAI221_X1 \mexu/_1154_ ( .A(\mexu/_0408_ ), .B1(\mexu/_0404_ ), .B2(\mexu/_0412_ ), .C1(\mexu/_0414_ ), .C2(\mexu/_0418_ ), .ZN(\mexu/_1010_ ) );
NAND2_X1 \mexu/_1155_ ( .A1(\mexu/_0175_ ), .A2(\mexu/_0174_ ), .ZN(\mexu/_0419_ ) );
OAI21_X1 \mexu/_1156_ ( .A(\mexu/_0419_ ), .B1(\mexu/_0414_ ), .B2(\mexu/_0417_ ), .ZN(\mexu/_0420_ ) );
BUF_X4 \mexu/_1157_ ( .A(\mexu/_0399_ ), .Z(\mexu/_0421_ ) );
NAND2_X1 \mexu/_1158_ ( .A1(\mexu/_0420_ ), .A2(\mexu/_0421_ ), .ZN(\mexu/_0422_ ) );
OAI21_X1 \mexu/_1159_ ( .A(\mexu/_0419_ ), .B1(\mexu/_0414_ ), .B2(\mexu/_0415_ ), .ZN(\mexu/_0423_ ) );
NAND2_X1 \mexu/_1160_ ( .A1(\mexu/_0423_ ), .A2(\mexu/_0400_ ), .ZN(\mexu/_0424_ ) );
BUF_X4 \mexu/_1161_ ( .A(\mexu/_0368_ ), .Z(\mexu/_0425_ ) );
NAND3_X1 \mexu/_1162_ ( .A1(\mexu/_0425_ ), .A2(\mexu/_0175_ ), .A3(\mexu/_0387_ ), .ZN(\mexu/_0426_ ) );
AND2_X1 \mexu/_1163_ ( .A1(\mexu/_0975_ ), .A2(\mexu/_0976_ ), .ZN(\mexu/_0427_ ) );
BUF_X4 \mexu/_1164_ ( .A(\mexu/_0427_ ), .Z(\mexu/_0428_ ) );
AND2_X1 \mexu/_1165_ ( .A1(\mexu/_0409_ ), .A2(\mexu/_0404_ ), .ZN(\mexu/_0429_ ) );
BUF_X4 \mexu/_1166_ ( .A(\mexu/_0429_ ), .Z(\mexu/_0430_ ) );
BUF_X4 \mexu/_1167_ ( .A(\mexu/_0430_ ), .Z(\mexu/_0431_ ) );
NAND4_X1 \mexu/_1168_ ( .A1(\mexu/_0425_ ), .A2(\mexu/_0977_ ), .A3(\mexu/_0428_ ), .A4(\mexu/_0431_ ), .ZN(\mexu/_0432_ ) );
NAND4_X1 \mexu/_1169_ ( .A1(\mexu/_0422_ ), .A2(\mexu/_0424_ ), .A3(\mexu/_0426_ ), .A4(\mexu/_0432_ ), .ZN(\mexu/_1011_ ) );
OAI221_X1 \mexu/_1170_ ( .A(\mexu/_0419_ ), .B1(\mexu/_0173_ ), .B2(\mexu/_0174_ ), .C1(\mexu/_0421_ ), .C2(\mexu/_0400_ ), .ZN(\mexu/_0433_ ) );
INV_X1 \mexu/_1171_ ( .A(\mexu/_0433_ ), .ZN(\mexu/_1012_ ) );
OAI21_X1 \mexu/_1172_ ( .A(\mexu/_0412_ ), .B1(\mexu/_0401_ ), .B2(\mexu/_0410_ ), .ZN(\mexu/_1013_ ) );
INV_X1 \mexu/_1173_ ( .A(\mexu/_0377_ ), .ZN(\mexu/_0434_ ) );
INV_X1 \mexu/_1174_ ( .A(\mexu/_0187_ ), .ZN(\mexu/_0435_ ) );
INV_X1 \mexu/_1175_ ( .A(\mexu/_0176_ ), .ZN(\mexu/_0436_ ) );
AOI21_X1 \mexu/_1176_ ( .A(\mexu/_0434_ ), .B1(\mexu/_0435_ ), .B2(\mexu/_0436_ ), .ZN(\mexu/_1014_ ) );
NOR4_X1 \mexu/_1177_ ( .A1(\mexu/_0175_ ), .A2(\mexu/_0173_ ), .A3(\mexu/_0174_ ), .A4(\mexu/_0187_ ), .ZN(\mexu/_1015_ ) );
NAND2_X1 \mexu/_1178_ ( .A1(\mexu/_0405_ ), .A2(\mexu/_0376_ ), .ZN(\mexu/_0437_ ) );
OAI21_X1 \mexu/_1179_ ( .A(\mexu/_0437_ ), .B1(\mexu/_0410_ ), .B2(\mexu/_0173_ ), .ZN(\mexu/_1016_ ) );
INV_X1 \mexu/_1180_ ( .A(\mexu/_0213_ ), .ZN(\mexu/_0438_ ) );
NAND4_X2 \mexu/_1181_ ( .A1(\mexu/_0379_ ), .A2(\mexu/_0438_ ), .A3(\mexu/_0395_ ), .A4(\mexu/_0384_ ), .ZN(\mexu/_0439_ ) );
NOR2_X1 \mexu/_1182_ ( .A1(\mexu/_0439_ ), .A2(\mexu/_0399_ ), .ZN(\mexu/_0440_ ) );
AOI221_X4 \mexu/_1183_ ( .A(\mexu/_0390_ ), .B1(\mexu/_0381_ ), .B2(\mexu/_0387_ ), .C1(\mexu/_0368_ ), .C2(\mexu/_0371_ ), .ZN(\mexu/_0441_ ) );
AND2_X1 \mexu/_1184_ ( .A1(\mexu/_0440_ ), .A2(\mexu/_0441_ ), .ZN(\mexu/_0442_ ) );
BUF_X4 \mexu/_1185_ ( .A(\mexu/_0442_ ), .Z(\mexu/_0443_ ) );
AND3_X1 \mexu/_1186_ ( .A1(\mexu/_0366_ ), .A2(\mexu/_0367_ ), .A3(\mexu/_0977_ ), .ZN(\mexu/_0444_ ) );
AND2_X1 \mexu/_1187_ ( .A1(\mexu/_0444_ ), .A2(\mexu/_0427_ ), .ZN(\mexu/_0445_ ) );
AND2_X1 \mexu/_1188_ ( .A1(\mexu/_0445_ ), .A2(\mexu/_0377_ ), .ZN(\mexu/_0446_ ) );
BUF_X4 \mexu/_1189_ ( .A(\mexu/_0446_ ), .Z(\mexu/_0447_ ) );
OAI21_X1 \mexu/_1190_ ( .A(\mexu/_1052_ ), .B1(\mexu/_0443_ ), .B2(\mexu/_0447_ ), .ZN(\mexu/_0448_ ) );
NAND4_X1 \mexu/_1191_ ( .A1(\mexu/_0425_ ), .A2(\mexu/_0140_ ), .A3(\mexu/_0372_ ), .A4(\mexu/_0431_ ), .ZN(\mexu/_0449_ ) );
BUF_X4 \mexu/_1192_ ( .A(\mexu/_0440_ ), .Z(\mexu/_0450_ ) );
OAI211_X2 \mexu/_1193_ ( .A(\mexu/_0448_ ), .B(\mexu/_0449_ ), .C1(\mexu/_0436_ ), .C2(\mexu/_0450_ ), .ZN(\mexu/_0108_ ) );
OAI21_X1 \mexu/_1194_ ( .A(\mexu/_1063_ ), .B1(\mexu/_0443_ ), .B2(\mexu/_0447_ ), .ZN(\mexu/_0451_ ) );
NAND4_X1 \mexu/_1195_ ( .A1(\mexu/_0425_ ), .A2(\mexu/_0151_ ), .A3(\mexu/_0372_ ), .A4(\mexu/_0430_ ), .ZN(\mexu/_0452_ ) );
OAI211_X2 \mexu/_1196_ ( .A(\mexu/_0451_ ), .B(\mexu/_0452_ ), .C1(\mexu/_0435_ ), .C2(\mexu/_0450_ ), .ZN(\mexu/_0119_ ) );
OAI21_X1 \mexu/_1197_ ( .A(\mexu/_1074_ ), .B1(\mexu/_0443_ ), .B2(\mexu/_0447_ ), .ZN(\mexu/_0453_ ) );
BUF_X4 \mexu/_1198_ ( .A(\mexu/_0391_ ), .Z(\mexu/_0454_ ) );
OAI21_X1 \mexu/_1199_ ( .A(\mexu/_0198_ ), .B1(\mexu/_0439_ ), .B2(\mexu/_0416_ ), .ZN(\mexu/_0455_ ) );
NAND4_X1 \mexu/_1200_ ( .A1(\mexu/_0425_ ), .A2(\mexu/_0162_ ), .A3(\mexu/_0372_ ), .A4(\mexu/_0431_ ), .ZN(\mexu/_0456_ ) );
NAND4_X1 \mexu/_1201_ ( .A1(\mexu/_0453_ ), .A2(\mexu/_0454_ ), .A3(\mexu/_0455_ ), .A4(\mexu/_0456_ ), .ZN(\mexu/_0130_ ) );
BUF_X4 \mexu/_1202_ ( .A(\mexu/_0442_ ), .Z(\mexu/_0457_ ) );
BUF_X4 \mexu/_1203_ ( .A(\mexu/_0446_ ), .Z(\mexu/_0458_ ) );
OAI21_X1 \mexu/_1204_ ( .A(\mexu/_1077_ ), .B1(\mexu/_0457_ ), .B2(\mexu/_0458_ ), .ZN(\mexu/_0459_ ) );
BUF_X4 \mexu/_1205_ ( .A(\mexu/_0439_ ), .Z(\mexu/_0460_ ) );
OAI21_X1 \mexu/_1206_ ( .A(\mexu/_0201_ ), .B1(\mexu/_0460_ ), .B2(\mexu/_0421_ ), .ZN(\mexu/_0461_ ) );
BUF_X4 \mexu/_1207_ ( .A(\mexu/_0430_ ), .Z(\mexu/_0462_ ) );
NAND4_X1 \mexu/_1208_ ( .A1(\mexu/_0373_ ), .A2(\mexu/_0165_ ), .A3(\mexu/_0374_ ), .A4(\mexu/_0462_ ), .ZN(\mexu/_0463_ ) );
NAND3_X1 \mexu/_1209_ ( .A1(\mexu/_0459_ ), .A2(\mexu/_0461_ ), .A3(\mexu/_0463_ ), .ZN(\mexu/_0133_ ) );
OAI21_X1 \mexu/_1210_ ( .A(\mexu/_1078_ ), .B1(\mexu/_0457_ ), .B2(\mexu/_0458_ ), .ZN(\mexu/_0464_ ) );
OAI21_X1 \mexu/_1211_ ( .A(\mexu/_0202_ ), .B1(\mexu/_0460_ ), .B2(\mexu/_0421_ ), .ZN(\mexu/_0465_ ) );
BUF_X4 \mexu/_1212_ ( .A(\mexu/_0444_ ), .Z(\mexu/_0466_ ) );
BUF_X4 \mexu/_1213_ ( .A(\mexu/_0466_ ), .Z(\mexu/_0467_ ) );
BUF_X4 \mexu/_1214_ ( .A(\mexu/_0427_ ), .Z(\mexu/_0468_ ) );
BUF_X4 \mexu/_1215_ ( .A(\mexu/_0468_ ), .Z(\mexu/_0469_ ) );
NAND4_X1 \mexu/_1216_ ( .A1(\mexu/_0467_ ), .A2(\mexu/_0166_ ), .A3(\mexu/_0469_ ), .A4(\mexu/_0462_ ), .ZN(\mexu/_0470_ ) );
NAND3_X1 \mexu/_1217_ ( .A1(\mexu/_0464_ ), .A2(\mexu/_0465_ ), .A3(\mexu/_0470_ ), .ZN(\mexu/_0134_ ) );
OAI21_X1 \mexu/_1218_ ( .A(\mexu/_1079_ ), .B1(\mexu/_0443_ ), .B2(\mexu/_0447_ ), .ZN(\mexu/_0471_ ) );
NAND4_X1 \mexu/_1219_ ( .A1(\mexu/_0466_ ), .A2(\mexu/_0167_ ), .A3(\mexu/_0468_ ), .A4(\mexu/_0430_ ), .ZN(\mexu/_0472_ ) );
OAI211_X2 \mexu/_1220_ ( .A(\mexu/_0471_ ), .B(\mexu/_0472_ ), .C1(\mexu/_0415_ ), .C2(\mexu/_0450_ ), .ZN(\mexu/_0135_ ) );
BUF_X4 \mexu/_1221_ ( .A(\mexu/_0441_ ), .Z(\mexu/_0473_ ) );
NAND3_X1 \mexu/_1222_ ( .A1(\mexu/_0450_ ), .A2(\mexu/_1080_ ), .A3(\mexu/_0473_ ), .ZN(\mexu/_0474_ ) );
BUF_X4 \mexu/_1223_ ( .A(\mexu/_0439_ ), .Z(\mexu/_0475_ ) );
BUF_X4 \mexu/_1224_ ( .A(\mexu/_0399_ ), .Z(\mexu/_0476_ ) );
OAI21_X1 \mexu/_1225_ ( .A(\mexu/_0204_ ), .B1(\mexu/_0475_ ), .B2(\mexu/_0476_ ), .ZN(\mexu/_0477_ ) );
BUF_X4 \mexu/_1226_ ( .A(\mexu/_0430_ ), .Z(\mexu/_0478_ ) );
NAND4_X1 \mexu/_1227_ ( .A1(\mexu/_0467_ ), .A2(\mexu/_0168_ ), .A3(\mexu/_0469_ ), .A4(\mexu/_0478_ ), .ZN(\mexu/_0479_ ) );
BUF_X4 \mexu/_1228_ ( .A(\mexu/_0466_ ), .Z(\mexu/_0480_ ) );
NAND4_X1 \mexu/_1229_ ( .A1(\mexu/_0480_ ), .A2(\mexu/_1080_ ), .A3(\mexu/_0428_ ), .A4(\mexu/_0378_ ), .ZN(\mexu/_0481_ ) );
NAND4_X1 \mexu/_1230_ ( .A1(\mexu/_0474_ ), .A2(\mexu/_0477_ ), .A3(\mexu/_0479_ ), .A4(\mexu/_0481_ ), .ZN(\mexu/_0136_ ) );
OAI21_X1 \mexu/_1231_ ( .A(\mexu/_1081_ ), .B1(\mexu/_0457_ ), .B2(\mexu/_0458_ ), .ZN(\mexu/_0482_ ) );
OAI21_X1 \mexu/_1232_ ( .A(\mexu/_0205_ ), .B1(\mexu/_0460_ ), .B2(\mexu/_0421_ ), .ZN(\mexu/_0483_ ) );
NAND4_X1 \mexu/_1233_ ( .A1(\mexu/_0467_ ), .A2(\mexu/_0169_ ), .A3(\mexu/_0469_ ), .A4(\mexu/_0462_ ), .ZN(\mexu/_0484_ ) );
NAND3_X1 \mexu/_1234_ ( .A1(\mexu/_0482_ ), .A2(\mexu/_0483_ ), .A3(\mexu/_0484_ ), .ZN(\mexu/_0137_ ) );
OAI21_X1 \mexu/_1235_ ( .A(\mexu/_1082_ ), .B1(\mexu/_0457_ ), .B2(\mexu/_0458_ ), .ZN(\mexu/_0485_ ) );
OAI21_X1 \mexu/_1236_ ( .A(\mexu/_0206_ ), .B1(\mexu/_0460_ ), .B2(\mexu/_0421_ ), .ZN(\mexu/_0486_ ) );
NAND4_X1 \mexu/_1237_ ( .A1(\mexu/_0373_ ), .A2(\mexu/_0170_ ), .A3(\mexu/_0374_ ), .A4(\mexu/_0462_ ), .ZN(\mexu/_0487_ ) );
NAND3_X1 \mexu/_1238_ ( .A1(\mexu/_0485_ ), .A2(\mexu/_0486_ ), .A3(\mexu/_0487_ ), .ZN(\mexu/_0138_ ) );
OAI21_X1 \mexu/_1239_ ( .A(\mexu/_1083_ ), .B1(\mexu/_0457_ ), .B2(\mexu/_0458_ ), .ZN(\mexu/_0488_ ) );
OAI21_X1 \mexu/_1240_ ( .A(\mexu/_0207_ ), .B1(\mexu/_0460_ ), .B2(\mexu/_0421_ ), .ZN(\mexu/_0489_ ) );
NAND4_X1 \mexu/_1241_ ( .A1(\mexu/_0373_ ), .A2(\mexu/_0171_ ), .A3(\mexu/_0374_ ), .A4(\mexu/_0462_ ), .ZN(\mexu/_0490_ ) );
NAND3_X1 \mexu/_1242_ ( .A1(\mexu/_0488_ ), .A2(\mexu/_0489_ ), .A3(\mexu/_0490_ ), .ZN(\mexu/_0139_ ) );
OAI21_X1 \mexu/_1243_ ( .A(\mexu/_1053_ ), .B1(\mexu/_0443_ ), .B2(\mexu/_0447_ ), .ZN(\mexu/_0491_ ) );
NAND4_X1 \mexu/_1244_ ( .A1(\mexu/_0425_ ), .A2(\mexu/_0141_ ), .A3(\mexu/_0372_ ), .A4(\mexu/_0430_ ), .ZN(\mexu/_0492_ ) );
OAI211_X2 \mexu/_1245_ ( .A(\mexu/_0491_ ), .B(\mexu/_0492_ ), .C1(\mexu/_0417_ ), .C2(\mexu/_0450_ ), .ZN(\mexu/_0109_ ) );
NAND3_X1 \mexu/_1246_ ( .A1(\mexu/_0450_ ), .A2(\mexu/_1054_ ), .A3(\mexu/_0473_ ), .ZN(\mexu/_0493_ ) );
OAI21_X1 \mexu/_1247_ ( .A(\mexu/_0178_ ), .B1(\mexu/_0475_ ), .B2(\mexu/_0476_ ), .ZN(\mexu/_0494_ ) );
NAND4_X1 \mexu/_1248_ ( .A1(\mexu/_0467_ ), .A2(\mexu/_0142_ ), .A3(\mexu/_0469_ ), .A4(\mexu/_0478_ ), .ZN(\mexu/_0495_ ) );
NAND4_X1 \mexu/_1249_ ( .A1(\mexu/_0480_ ), .A2(\mexu/_1054_ ), .A3(\mexu/_0428_ ), .A4(\mexu/_0378_ ), .ZN(\mexu/_0496_ ) );
NAND4_X1 \mexu/_1250_ ( .A1(\mexu/_0493_ ), .A2(\mexu/_0494_ ), .A3(\mexu/_0495_ ), .A4(\mexu/_0496_ ), .ZN(\mexu/_0110_ ) );
OAI21_X1 \mexu/_1251_ ( .A(\mexu/_1055_ ), .B1(\mexu/_0457_ ), .B2(\mexu/_0458_ ), .ZN(\mexu/_0497_ ) );
OAI21_X1 \mexu/_1252_ ( .A(\mexu/_0179_ ), .B1(\mexu/_0460_ ), .B2(\mexu/_0421_ ), .ZN(\mexu/_0498_ ) );
NAND4_X1 \mexu/_1253_ ( .A1(\mexu/_0467_ ), .A2(\mexu/_0143_ ), .A3(\mexu/_0469_ ), .A4(\mexu/_0462_ ), .ZN(\mexu/_0499_ ) );
NAND3_X1 \mexu/_1254_ ( .A1(\mexu/_0497_ ), .A2(\mexu/_0498_ ), .A3(\mexu/_0499_ ), .ZN(\mexu/_0111_ ) );
OAI21_X1 \mexu/_1255_ ( .A(\mexu/_1056_ ), .B1(\mexu/_0457_ ), .B2(\mexu/_0458_ ), .ZN(\mexu/_0500_ ) );
OAI21_X1 \mexu/_1256_ ( .A(\mexu/_0180_ ), .B1(\mexu/_0460_ ), .B2(\mexu/_0421_ ), .ZN(\mexu/_0501_ ) );
NAND4_X1 \mexu/_1257_ ( .A1(\mexu/_0373_ ), .A2(\mexu/_0144_ ), .A3(\mexu/_0374_ ), .A4(\mexu/_0462_ ), .ZN(\mexu/_0502_ ) );
NAND3_X1 \mexu/_1258_ ( .A1(\mexu/_0500_ ), .A2(\mexu/_0501_ ), .A3(\mexu/_0502_ ), .ZN(\mexu/_0112_ ) );
NAND3_X1 \mexu/_1259_ ( .A1(\mexu/_0450_ ), .A2(\mexu/_1057_ ), .A3(\mexu/_0473_ ), .ZN(\mexu/_0503_ ) );
OAI21_X1 \mexu/_1260_ ( .A(\mexu/_0181_ ), .B1(\mexu/_0475_ ), .B2(\mexu/_0416_ ), .ZN(\mexu/_0504_ ) );
NAND4_X1 \mexu/_1261_ ( .A1(\mexu/_0467_ ), .A2(\mexu/_0145_ ), .A3(\mexu/_0469_ ), .A4(\mexu/_0478_ ), .ZN(\mexu/_0505_ ) );
NAND4_X1 \mexu/_1262_ ( .A1(\mexu/_0480_ ), .A2(\mexu/_1057_ ), .A3(\mexu/_0428_ ), .A4(\mexu/_0378_ ), .ZN(\mexu/_0506_ ) );
NAND4_X1 \mexu/_1263_ ( .A1(\mexu/_0503_ ), .A2(\mexu/_0504_ ), .A3(\mexu/_0505_ ), .A4(\mexu/_0506_ ), .ZN(\mexu/_0113_ ) );
OAI21_X1 \mexu/_1264_ ( .A(\mexu/_1058_ ), .B1(\mexu/_0443_ ), .B2(\mexu/_0447_ ), .ZN(\mexu/_0507_ ) );
NAND4_X1 \mexu/_1265_ ( .A1(\mexu/_0425_ ), .A2(\mexu/_0146_ ), .A3(\mexu/_0372_ ), .A4(\mexu/_0430_ ), .ZN(\mexu/_0508_ ) );
INV_X1 \mexu/_1266_ ( .A(\mexu/_0182_ ), .ZN(\mexu/_0509_ ) );
OAI211_X2 \mexu/_1267_ ( .A(\mexu/_0507_ ), .B(\mexu/_0508_ ), .C1(\mexu/_0509_ ), .C2(\mexu/_0450_ ), .ZN(\mexu/_0114_ ) );
NAND3_X1 \mexu/_1268_ ( .A1(\mexu/_0450_ ), .A2(\mexu/_1059_ ), .A3(\mexu/_0473_ ), .ZN(\mexu/_0510_ ) );
OAI21_X1 \mexu/_1269_ ( .A(\mexu/_0183_ ), .B1(\mexu/_0475_ ), .B2(\mexu/_0416_ ), .ZN(\mexu/_0511_ ) );
NAND4_X1 \mexu/_1270_ ( .A1(\mexu/_0467_ ), .A2(\mexu/_0147_ ), .A3(\mexu/_0469_ ), .A4(\mexu/_0478_ ), .ZN(\mexu/_0512_ ) );
NAND4_X1 \mexu/_1271_ ( .A1(\mexu/_0480_ ), .A2(\mexu/_1059_ ), .A3(\mexu/_0428_ ), .A4(\mexu/_0378_ ), .ZN(\mexu/_0513_ ) );
NAND4_X1 \mexu/_1272_ ( .A1(\mexu/_0510_ ), .A2(\mexu/_0511_ ), .A3(\mexu/_0512_ ), .A4(\mexu/_0513_ ), .ZN(\mexu/_0115_ ) );
NAND3_X1 \mexu/_1273_ ( .A1(\mexu/_0450_ ), .A2(\mexu/_1060_ ), .A3(\mexu/_0473_ ), .ZN(\mexu/_0514_ ) );
OAI21_X1 \mexu/_1274_ ( .A(\mexu/_0184_ ), .B1(\mexu/_0439_ ), .B2(\mexu/_0416_ ), .ZN(\mexu/_0515_ ) );
NAND4_X1 \mexu/_1275_ ( .A1(\mexu/_0467_ ), .A2(\mexu/_0148_ ), .A3(\mexu/_0469_ ), .A4(\mexu/_0478_ ), .ZN(\mexu/_0516_ ) );
NAND4_X1 \mexu/_1276_ ( .A1(\mexu/_0480_ ), .A2(\mexu/_1060_ ), .A3(\mexu/_0468_ ), .A4(\mexu/_0378_ ), .ZN(\mexu/_0517_ ) );
NAND4_X1 \mexu/_1277_ ( .A1(\mexu/_0514_ ), .A2(\mexu/_0515_ ), .A3(\mexu/_0516_ ), .A4(\mexu/_0517_ ), .ZN(\mexu/_0116_ ) );
OAI21_X1 \mexu/_1278_ ( .A(\mexu/_1061_ ), .B1(\mexu/_0457_ ), .B2(\mexu/_0458_ ), .ZN(\mexu/_0518_ ) );
OAI21_X1 \mexu/_1279_ ( .A(\mexu/_0185_ ), .B1(\mexu/_0460_ ), .B2(\mexu/_0421_ ), .ZN(\mexu/_0519_ ) );
NAND4_X1 \mexu/_1280_ ( .A1(\mexu/_0373_ ), .A2(\mexu/_0149_ ), .A3(\mexu/_0374_ ), .A4(\mexu/_0462_ ), .ZN(\mexu/_0520_ ) );
NAND3_X1 \mexu/_1281_ ( .A1(\mexu/_0518_ ), .A2(\mexu/_0519_ ), .A3(\mexu/_0520_ ), .ZN(\mexu/_0117_ ) );
OAI21_X1 \mexu/_1282_ ( .A(\mexu/_1062_ ), .B1(\mexu/_0457_ ), .B2(\mexu/_0458_ ), .ZN(\mexu/_0521_ ) );
OAI21_X1 \mexu/_1283_ ( .A(\mexu/_0186_ ), .B1(\mexu/_0460_ ), .B2(\mexu/_0476_ ), .ZN(\mexu/_0522_ ) );
NAND4_X1 \mexu/_1284_ ( .A1(\mexu/_0373_ ), .A2(\mexu/_0150_ ), .A3(\mexu/_0374_ ), .A4(\mexu/_0462_ ), .ZN(\mexu/_0523_ ) );
NAND3_X1 \mexu/_1285_ ( .A1(\mexu/_0521_ ), .A2(\mexu/_0522_ ), .A3(\mexu/_0523_ ), .ZN(\mexu/_0118_ ) );
NAND3_X1 \mexu/_1286_ ( .A1(\mexu/_0440_ ), .A2(\mexu/_1064_ ), .A3(\mexu/_0473_ ), .ZN(\mexu/_0524_ ) );
OAI21_X1 \mexu/_1287_ ( .A(\mexu/_0188_ ), .B1(\mexu/_0439_ ), .B2(\mexu/_0416_ ), .ZN(\mexu/_0525_ ) );
NAND4_X1 \mexu/_1288_ ( .A1(\mexu/_0467_ ), .A2(\mexu/_0152_ ), .A3(\mexu/_0469_ ), .A4(\mexu/_0431_ ), .ZN(\mexu/_0526_ ) );
NAND4_X1 \mexu/_1289_ ( .A1(\mexu/_0466_ ), .A2(\mexu/_1064_ ), .A3(\mexu/_0468_ ), .A4(\mexu/_0378_ ), .ZN(\mexu/_0527_ ) );
NAND4_X1 \mexu/_1290_ ( .A1(\mexu/_0524_ ), .A2(\mexu/_0525_ ), .A3(\mexu/_0526_ ), .A4(\mexu/_0527_ ), .ZN(\mexu/_0120_ ) );
NAND3_X1 \mexu/_1291_ ( .A1(\mexu/_0440_ ), .A2(\mexu/_1065_ ), .A3(\mexu/_0473_ ), .ZN(\mexu/_0528_ ) );
OAI21_X1 \mexu/_1292_ ( .A(\mexu/_0189_ ), .B1(\mexu/_0439_ ), .B2(\mexu/_0416_ ), .ZN(\mexu/_0529_ ) );
NAND4_X1 \mexu/_1293_ ( .A1(\mexu/_0467_ ), .A2(\mexu/_0153_ ), .A3(\mexu/_0469_ ), .A4(\mexu/_0431_ ), .ZN(\mexu/_0530_ ) );
NAND4_X1 \mexu/_1294_ ( .A1(\mexu/_0466_ ), .A2(\mexu/_1065_ ), .A3(\mexu/_0468_ ), .A4(\mexu/_0378_ ), .ZN(\mexu/_0531_ ) );
NAND4_X1 \mexu/_1295_ ( .A1(\mexu/_0528_ ), .A2(\mexu/_0529_ ), .A3(\mexu/_0530_ ), .A4(\mexu/_0531_ ), .ZN(\mexu/_0121_ ) );
OAI21_X1 \mexu/_1296_ ( .A(\mexu/_1066_ ), .B1(\mexu/_0457_ ), .B2(\mexu/_0458_ ), .ZN(\mexu/_0532_ ) );
OAI21_X1 \mexu/_1297_ ( .A(\mexu/_0190_ ), .B1(\mexu/_0460_ ), .B2(\mexu/_0476_ ), .ZN(\mexu/_0533_ ) );
NAND4_X1 \mexu/_1298_ ( .A1(\mexu/_0373_ ), .A2(\mexu/_0154_ ), .A3(\mexu/_0374_ ), .A4(\mexu/_0478_ ), .ZN(\mexu/_0534_ ) );
NAND3_X1 \mexu/_1299_ ( .A1(\mexu/_0532_ ), .A2(\mexu/_0533_ ), .A3(\mexu/_0534_ ), .ZN(\mexu/_0122_ ) );
NAND3_X1 \mexu/_1300_ ( .A1(\mexu/_0440_ ), .A2(\mexu/_1067_ ), .A3(\mexu/_0473_ ), .ZN(\mexu/_0535_ ) );
OAI21_X1 \mexu/_1301_ ( .A(\mexu/_0191_ ), .B1(\mexu/_0439_ ), .B2(\mexu/_0416_ ), .ZN(\mexu/_0536_ ) );
NAND4_X1 \mexu/_1302_ ( .A1(\mexu/_0480_ ), .A2(\mexu/_0155_ ), .A3(\mexu/_0428_ ), .A4(\mexu/_0431_ ), .ZN(\mexu/_0537_ ) );
NAND4_X1 \mexu/_1303_ ( .A1(\mexu/_0466_ ), .A2(\mexu/_1067_ ), .A3(\mexu/_0468_ ), .A4(\mexu/_0378_ ), .ZN(\mexu/_0538_ ) );
NAND4_X1 \mexu/_1304_ ( .A1(\mexu/_0535_ ), .A2(\mexu/_0536_ ), .A3(\mexu/_0537_ ), .A4(\mexu/_0538_ ), .ZN(\mexu/_0123_ ) );
NAND3_X1 \mexu/_1305_ ( .A1(\mexu/_0440_ ), .A2(\mexu/_1068_ ), .A3(\mexu/_0473_ ), .ZN(\mexu/_0539_ ) );
OAI21_X1 \mexu/_1306_ ( .A(\mexu/_0192_ ), .B1(\mexu/_0439_ ), .B2(\mexu/_0416_ ), .ZN(\mexu/_0540_ ) );
NAND4_X1 \mexu/_1307_ ( .A1(\mexu/_0480_ ), .A2(\mexu/_0156_ ), .A3(\mexu/_0428_ ), .A4(\mexu/_0431_ ), .ZN(\mexu/_0541_ ) );
NAND4_X1 \mexu/_1308_ ( .A1(\mexu/_0466_ ), .A2(\mexu/_1068_ ), .A3(\mexu/_0468_ ), .A4(\mexu/_0377_ ), .ZN(\mexu/_0542_ ) );
NAND4_X1 \mexu/_1309_ ( .A1(\mexu/_0539_ ), .A2(\mexu/_0540_ ), .A3(\mexu/_0541_ ), .A4(\mexu/_0542_ ), .ZN(\mexu/_0124_ ) );
OAI21_X1 \mexu/_1310_ ( .A(\mexu/_1069_ ), .B1(\mexu/_0443_ ), .B2(\mexu/_0447_ ), .ZN(\mexu/_0543_ ) );
OAI21_X1 \mexu/_1311_ ( .A(\mexu/_0193_ ), .B1(\mexu/_0475_ ), .B2(\mexu/_0476_ ), .ZN(\mexu/_0544_ ) );
NAND4_X1 \mexu/_1312_ ( .A1(\mexu/_0373_ ), .A2(\mexu/_0157_ ), .A3(\mexu/_0374_ ), .A4(\mexu/_0478_ ), .ZN(\mexu/_0545_ ) );
NAND3_X1 \mexu/_1313_ ( .A1(\mexu/_0543_ ), .A2(\mexu/_0544_ ), .A3(\mexu/_0545_ ), .ZN(\mexu/_0125_ ) );
OAI21_X1 \mexu/_1314_ ( .A(\mexu/_1070_ ), .B1(\mexu/_0443_ ), .B2(\mexu/_0447_ ), .ZN(\mexu/_0546_ ) );
OAI21_X1 \mexu/_1315_ ( .A(\mexu/_0194_ ), .B1(\mexu/_0475_ ), .B2(\mexu/_0476_ ), .ZN(\mexu/_0547_ ) );
NAND4_X1 \mexu/_1316_ ( .A1(\mexu/_0425_ ), .A2(\mexu/_0158_ ), .A3(\mexu/_0372_ ), .A4(\mexu/_0478_ ), .ZN(\mexu/_0548_ ) );
NAND3_X1 \mexu/_1317_ ( .A1(\mexu/_0546_ ), .A2(\mexu/_0547_ ), .A3(\mexu/_0548_ ), .ZN(\mexu/_0126_ ) );
NAND3_X1 \mexu/_1318_ ( .A1(\mexu/_0440_ ), .A2(\mexu/_1071_ ), .A3(\mexu/_0473_ ), .ZN(\mexu/_0549_ ) );
OAI21_X1 \mexu/_1319_ ( .A(\mexu/_0195_ ), .B1(\mexu/_0439_ ), .B2(\mexu/_0416_ ), .ZN(\mexu/_0550_ ) );
NAND4_X1 \mexu/_1320_ ( .A1(\mexu/_0480_ ), .A2(\mexu/_0159_ ), .A3(\mexu/_0428_ ), .A4(\mexu/_0431_ ), .ZN(\mexu/_0551_ ) );
NAND4_X1 \mexu/_1321_ ( .A1(\mexu/_0466_ ), .A2(\mexu/_1071_ ), .A3(\mexu/_0468_ ), .A4(\mexu/_0377_ ), .ZN(\mexu/_0552_ ) );
NAND4_X1 \mexu/_1322_ ( .A1(\mexu/_0549_ ), .A2(\mexu/_0550_ ), .A3(\mexu/_0551_ ), .A4(\mexu/_0552_ ), .ZN(\mexu/_0127_ ) );
OAI21_X1 \mexu/_1323_ ( .A(\mexu/_1072_ ), .B1(\mexu/_0443_ ), .B2(\mexu/_0447_ ), .ZN(\mexu/_0553_ ) );
OAI21_X1 \mexu/_1324_ ( .A(\mexu/_0196_ ), .B1(\mexu/_0475_ ), .B2(\mexu/_0476_ ), .ZN(\mexu/_0554_ ) );
NAND4_X1 \mexu/_1325_ ( .A1(\mexu/_0425_ ), .A2(\mexu/_0160_ ), .A3(\mexu/_0372_ ), .A4(\mexu/_0478_ ), .ZN(\mexu/_0555_ ) );
NAND3_X1 \mexu/_1326_ ( .A1(\mexu/_0553_ ), .A2(\mexu/_0554_ ), .A3(\mexu/_0555_ ), .ZN(\mexu/_0128_ ) );
OAI21_X1 \mexu/_1327_ ( .A(\mexu/_0197_ ), .B1(\mexu/_0475_ ), .B2(\mexu/_0476_ ), .ZN(\mexu/_0556_ ) );
NOR2_X1 \mexu/_1328_ ( .A1(\mexu/_0213_ ), .A2(\mexu/_0398_ ), .ZN(\mexu/_0557_ ) );
NAND4_X1 \mexu/_1329_ ( .A1(\mexu/_0385_ ), .A2(\mexu/_1073_ ), .A3(\mexu/_0557_ ), .A4(\mexu/_0441_ ), .ZN(\mexu/_0558_ ) );
NAND4_X1 \mexu/_1330_ ( .A1(\mexu/_0480_ ), .A2(\mexu/_0161_ ), .A3(\mexu/_0428_ ), .A4(\mexu/_0431_ ), .ZN(\mexu/_0559_ ) );
NAND4_X1 \mexu/_1331_ ( .A1(\mexu/_0466_ ), .A2(\mexu/_1073_ ), .A3(\mexu/_0468_ ), .A4(\mexu/_0377_ ), .ZN(\mexu/_0560_ ) );
NAND4_X1 \mexu/_1332_ ( .A1(\mexu/_0556_ ), .A2(\mexu/_0558_ ), .A3(\mexu/_0559_ ), .A4(\mexu/_0560_ ), .ZN(\mexu/_0129_ ) );
OAI21_X1 \mexu/_1333_ ( .A(\mexu/_0199_ ), .B1(\mexu/_0475_ ), .B2(\mexu/_0476_ ), .ZN(\mexu/_0561_ ) );
NAND4_X1 \mexu/_1334_ ( .A1(\mexu/_0385_ ), .A2(\mexu/_1075_ ), .A3(\mexu/_0557_ ), .A4(\mexu/_0441_ ), .ZN(\mexu/_0562_ ) );
NAND4_X1 \mexu/_1335_ ( .A1(\mexu/_0480_ ), .A2(\mexu/_0163_ ), .A3(\mexu/_0428_ ), .A4(\mexu/_0431_ ), .ZN(\mexu/_0563_ ) );
NAND4_X1 \mexu/_1336_ ( .A1(\mexu/_0466_ ), .A2(\mexu/_1075_ ), .A3(\mexu/_0468_ ), .A4(\mexu/_0377_ ), .ZN(\mexu/_0564_ ) );
NAND4_X1 \mexu/_1337_ ( .A1(\mexu/_0561_ ), .A2(\mexu/_0562_ ), .A3(\mexu/_0563_ ), .A4(\mexu/_0564_ ), .ZN(\mexu/_0131_ ) );
OAI21_X1 \mexu/_1338_ ( .A(\mexu/_1076_ ), .B1(\mexu/_0443_ ), .B2(\mexu/_0447_ ), .ZN(\mexu/_0565_ ) );
OAI21_X1 \mexu/_1339_ ( .A(\mexu/_0200_ ), .B1(\mexu/_0475_ ), .B2(\mexu/_0476_ ), .ZN(\mexu/_0566_ ) );
NAND4_X1 \mexu/_1340_ ( .A1(\mexu/_0425_ ), .A2(\mexu/_0164_ ), .A3(\mexu/_0372_ ), .A4(\mexu/_0478_ ), .ZN(\mexu/_0567_ ) );
NAND3_X1 \mexu/_1341_ ( .A1(\mexu/_0565_ ), .A2(\mexu/_0566_ ), .A3(\mexu/_0567_ ), .ZN(\mexu/_0132_ ) );
INV_X1 \mexu/_1342_ ( .A(\mexu/_0391_ ), .ZN(\mexu/_0568_ ) );
BUF_X4 \mexu/_1343_ ( .A(\mexu/_0568_ ), .Z(\mexu/_0569_ ) );
BUF_X4 \mexu/_1344_ ( .A(\mexu/_0394_ ), .Z(\mexu/_0570_ ) );
OAI21_X1 \mexu/_1345_ ( .A(\mexu/_0978_ ), .B1(\mexu/_0569_ ), .B2(\mexu/_0570_ ), .ZN(\mexu/_0571_ ) );
BUF_X4 \mexu/_1346_ ( .A(\mexu/_0395_ ), .Z(\mexu/_0572_ ) );
BUF_X4 \mexu/_1347_ ( .A(\mexu/_0384_ ), .Z(\mexu/_0573_ ) );
NAND4_X1 \mexu/_1348_ ( .A1(\mexu/_0454_ ), .A2(\mexu/_1020_ ), .A3(\mexu/_0572_ ), .A4(\mexu/_0573_ ), .ZN(\mexu/_0574_ ) );
NAND2_X1 \mexu/_1349_ ( .A1(\mexu/_0571_ ), .A2(\mexu/_0574_ ), .ZN(\mexu/_0076_ ) );
OAI21_X1 \mexu/_1350_ ( .A(\mexu/_0989_ ), .B1(\mexu/_0569_ ), .B2(\mexu/_0570_ ), .ZN(\mexu/_0575_ ) );
NAND4_X1 \mexu/_1351_ ( .A1(\mexu/_0454_ ), .A2(\mexu/_1031_ ), .A3(\mexu/_0572_ ), .A4(\mexu/_0573_ ), .ZN(\mexu/_0576_ ) );
NAND2_X1 \mexu/_1352_ ( .A1(\mexu/_0575_ ), .A2(\mexu/_0576_ ), .ZN(\mexu/_0087_ ) );
OAI21_X1 \mexu/_1353_ ( .A(\mexu/_1000_ ), .B1(\mexu/_0569_ ), .B2(\mexu/_0570_ ), .ZN(\mexu/_0577_ ) );
NAND4_X1 \mexu/_1354_ ( .A1(\mexu/_0454_ ), .A2(\mexu/_1042_ ), .A3(\mexu/_0572_ ), .A4(\mexu/_0573_ ), .ZN(\mexu/_0578_ ) );
NAND2_X1 \mexu/_1355_ ( .A1(\mexu/_0577_ ), .A2(\mexu/_0578_ ), .ZN(\mexu/_0098_ ) );
OAI21_X1 \mexu/_1356_ ( .A(\mexu/_1003_ ), .B1(\mexu/_0569_ ), .B2(\mexu/_0570_ ), .ZN(\mexu/_0579_ ) );
NAND4_X1 \mexu/_1357_ ( .A1(\mexu/_0454_ ), .A2(\mexu/_1045_ ), .A3(\mexu/_0572_ ), .A4(\mexu/_0573_ ), .ZN(\mexu/_0580_ ) );
NAND2_X1 \mexu/_1358_ ( .A1(\mexu/_0579_ ), .A2(\mexu/_0580_ ), .ZN(\mexu/_0101_ ) );
OAI21_X1 \mexu/_1359_ ( .A(\mexu/_1004_ ), .B1(\mexu/_0569_ ), .B2(\mexu/_0570_ ), .ZN(\mexu/_0581_ ) );
NAND4_X1 \mexu/_1360_ ( .A1(\mexu/_0454_ ), .A2(\mexu/_1046_ ), .A3(\mexu/_0572_ ), .A4(\mexu/_0573_ ), .ZN(\mexu/_0582_ ) );
NAND2_X1 \mexu/_1361_ ( .A1(\mexu/_0581_ ), .A2(\mexu/_0582_ ), .ZN(\mexu/_0102_ ) );
OAI21_X1 \mexu/_1362_ ( .A(\mexu/_1005_ ), .B1(\mexu/_0569_ ), .B2(\mexu/_0570_ ), .ZN(\mexu/_0583_ ) );
NAND4_X1 \mexu/_1363_ ( .A1(\mexu/_0454_ ), .A2(\mexu/_1047_ ), .A3(\mexu/_0572_ ), .A4(\mexu/_0573_ ), .ZN(\mexu/_0584_ ) );
NAND2_X1 \mexu/_1364_ ( .A1(\mexu/_0583_ ), .A2(\mexu/_0584_ ), .ZN(\mexu/_0103_ ) );
OAI21_X1 \mexu/_1365_ ( .A(\mexu/_1006_ ), .B1(\mexu/_0569_ ), .B2(\mexu/_0570_ ), .ZN(\mexu/_0585_ ) );
NAND4_X1 \mexu/_1366_ ( .A1(\mexu/_0454_ ), .A2(\mexu/_1048_ ), .A3(\mexu/_0572_ ), .A4(\mexu/_0573_ ), .ZN(\mexu/_0586_ ) );
NAND2_X1 \mexu/_1367_ ( .A1(\mexu/_0585_ ), .A2(\mexu/_0586_ ), .ZN(\mexu/_0104_ ) );
OAI21_X1 \mexu/_1368_ ( .A(\mexu/_1007_ ), .B1(\mexu/_0569_ ), .B2(\mexu/_0570_ ), .ZN(\mexu/_0587_ ) );
NAND4_X1 \mexu/_1369_ ( .A1(\mexu/_0454_ ), .A2(\mexu/_1049_ ), .A3(\mexu/_0572_ ), .A4(\mexu/_0573_ ), .ZN(\mexu/_0588_ ) );
NAND2_X1 \mexu/_1370_ ( .A1(\mexu/_0587_ ), .A2(\mexu/_0588_ ), .ZN(\mexu/_0105_ ) );
OAI21_X1 \mexu/_1371_ ( .A(\mexu/_1008_ ), .B1(\mexu/_0569_ ), .B2(\mexu/_0570_ ), .ZN(\mexu/_0589_ ) );
BUF_X4 \mexu/_1372_ ( .A(\mexu/_0391_ ), .Z(\mexu/_0590_ ) );
NAND4_X1 \mexu/_1373_ ( .A1(\mexu/_0590_ ), .A2(\mexu/_1050_ ), .A3(\mexu/_0572_ ), .A4(\mexu/_0573_ ), .ZN(\mexu/_0591_ ) );
NAND2_X1 \mexu/_1374_ ( .A1(\mexu/_0589_ ), .A2(\mexu/_0591_ ), .ZN(\mexu/_0106_ ) );
OAI21_X1 \mexu/_1375_ ( .A(\mexu/_1009_ ), .B1(\mexu/_0569_ ), .B2(\mexu/_0570_ ), .ZN(\mexu/_0592_ ) );
BUF_X4 \mexu/_1376_ ( .A(\mexu/_0384_ ), .Z(\mexu/_0593_ ) );
NAND4_X1 \mexu/_1377_ ( .A1(\mexu/_0590_ ), .A2(\mexu/_1051_ ), .A3(\mexu/_0572_ ), .A4(\mexu/_0593_ ), .ZN(\mexu/_0594_ ) );
NAND2_X1 \mexu/_1378_ ( .A1(\mexu/_0592_ ), .A2(\mexu/_0594_ ), .ZN(\mexu/_0107_ ) );
BUF_X4 \mexu/_1379_ ( .A(\mexu/_0568_ ), .Z(\mexu/_0595_ ) );
BUF_X4 \mexu/_1380_ ( .A(\mexu/_0394_ ), .Z(\mexu/_0596_ ) );
OAI21_X1 \mexu/_1381_ ( .A(\mexu/_0979_ ), .B1(\mexu/_0595_ ), .B2(\mexu/_0596_ ), .ZN(\mexu/_0597_ ) );
BUF_X4 \mexu/_1382_ ( .A(\mexu/_0395_ ), .Z(\mexu/_0598_ ) );
NAND4_X1 \mexu/_1383_ ( .A1(\mexu/_0590_ ), .A2(\mexu/_1021_ ), .A3(\mexu/_0598_ ), .A4(\mexu/_0593_ ), .ZN(\mexu/_0599_ ) );
NAND2_X1 \mexu/_1384_ ( .A1(\mexu/_0597_ ), .A2(\mexu/_0599_ ), .ZN(\mexu/_0077_ ) );
OAI21_X1 \mexu/_1385_ ( .A(\mexu/_0980_ ), .B1(\mexu/_0595_ ), .B2(\mexu/_0596_ ), .ZN(\mexu/_0600_ ) );
NAND4_X1 \mexu/_1386_ ( .A1(\mexu/_0590_ ), .A2(\mexu/_1022_ ), .A3(\mexu/_0598_ ), .A4(\mexu/_0593_ ), .ZN(\mexu/_0601_ ) );
NAND2_X1 \mexu/_1387_ ( .A1(\mexu/_0600_ ), .A2(\mexu/_0601_ ), .ZN(\mexu/_0078_ ) );
OAI21_X1 \mexu/_1388_ ( .A(\mexu/_0981_ ), .B1(\mexu/_0595_ ), .B2(\mexu/_0596_ ), .ZN(\mexu/_0602_ ) );
NAND4_X1 \mexu/_1389_ ( .A1(\mexu/_0590_ ), .A2(\mexu/_1023_ ), .A3(\mexu/_0598_ ), .A4(\mexu/_0593_ ), .ZN(\mexu/_0603_ ) );
NAND2_X1 \mexu/_1390_ ( .A1(\mexu/_0602_ ), .A2(\mexu/_0603_ ), .ZN(\mexu/_0079_ ) );
OAI21_X1 \mexu/_1391_ ( .A(\mexu/_0982_ ), .B1(\mexu/_0595_ ), .B2(\mexu/_0596_ ), .ZN(\mexu/_0604_ ) );
NAND4_X1 \mexu/_1392_ ( .A1(\mexu/_0590_ ), .A2(\mexu/_1024_ ), .A3(\mexu/_0598_ ), .A4(\mexu/_0593_ ), .ZN(\mexu/_0605_ ) );
NAND2_X1 \mexu/_1393_ ( .A1(\mexu/_0604_ ), .A2(\mexu/_0605_ ), .ZN(\mexu/_0080_ ) );
OAI21_X1 \mexu/_1394_ ( .A(\mexu/_0983_ ), .B1(\mexu/_0595_ ), .B2(\mexu/_0596_ ), .ZN(\mexu/_0606_ ) );
NAND4_X1 \mexu/_1395_ ( .A1(\mexu/_0590_ ), .A2(\mexu/_1025_ ), .A3(\mexu/_0598_ ), .A4(\mexu/_0593_ ), .ZN(\mexu/_0607_ ) );
NAND2_X1 \mexu/_1396_ ( .A1(\mexu/_0606_ ), .A2(\mexu/_0607_ ), .ZN(\mexu/_0081_ ) );
OAI21_X1 \mexu/_1397_ ( .A(\mexu/_0984_ ), .B1(\mexu/_0568_ ), .B2(\mexu/_0394_ ), .ZN(\mexu/_0608_ ) );
NAND2_X1 \mexu/_1398_ ( .A1(\mexu/_0396_ ), .A2(\mexu/_0573_ ), .ZN(\mexu/_0609_ ) );
INV_X1 \mexu/_1399_ ( .A(\mexu/_1026_ ), .ZN(\mexu/_0610_ ) );
OAI21_X1 \mexu/_1400_ ( .A(\mexu/_0608_ ), .B1(\mexu/_0609_ ), .B2(\mexu/_0610_ ), .ZN(\mexu/_0082_ ) );
OAI21_X1 \mexu/_1401_ ( .A(\mexu/_0985_ ), .B1(\mexu/_0595_ ), .B2(\mexu/_0596_ ), .ZN(\mexu/_0611_ ) );
NAND4_X1 \mexu/_1402_ ( .A1(\mexu/_0590_ ), .A2(\mexu/_1027_ ), .A3(\mexu/_0598_ ), .A4(\mexu/_0593_ ), .ZN(\mexu/_0612_ ) );
NAND2_X1 \mexu/_1403_ ( .A1(\mexu/_0611_ ), .A2(\mexu/_0612_ ), .ZN(\mexu/_0083_ ) );
OAI21_X1 \mexu/_1404_ ( .A(\mexu/_0986_ ), .B1(\mexu/_0595_ ), .B2(\mexu/_0596_ ), .ZN(\mexu/_0613_ ) );
NAND4_X1 \mexu/_1405_ ( .A1(\mexu/_0590_ ), .A2(\mexu/_1028_ ), .A3(\mexu/_0598_ ), .A4(\mexu/_0593_ ), .ZN(\mexu/_0614_ ) );
NAND2_X1 \mexu/_1406_ ( .A1(\mexu/_0613_ ), .A2(\mexu/_0614_ ), .ZN(\mexu/_0084_ ) );
OAI21_X1 \mexu/_1407_ ( .A(\mexu/_0987_ ), .B1(\mexu/_0595_ ), .B2(\mexu/_0596_ ), .ZN(\mexu/_0615_ ) );
NAND4_X1 \mexu/_1408_ ( .A1(\mexu/_0590_ ), .A2(\mexu/_1029_ ), .A3(\mexu/_0598_ ), .A4(\mexu/_0593_ ), .ZN(\mexu/_0616_ ) );
NAND2_X1 \mexu/_1409_ ( .A1(\mexu/_0615_ ), .A2(\mexu/_0616_ ), .ZN(\mexu/_0085_ ) );
OAI21_X1 \mexu/_1410_ ( .A(\mexu/_0988_ ), .B1(\mexu/_0595_ ), .B2(\mexu/_0596_ ), .ZN(\mexu/_0617_ ) );
BUF_X4 \mexu/_1411_ ( .A(\mexu/_0391_ ), .Z(\mexu/_0618_ ) );
NAND4_X1 \mexu/_1412_ ( .A1(\mexu/_0618_ ), .A2(\mexu/_1030_ ), .A3(\mexu/_0598_ ), .A4(\mexu/_0593_ ), .ZN(\mexu/_0619_ ) );
NAND2_X1 \mexu/_1413_ ( .A1(\mexu/_0617_ ), .A2(\mexu/_0619_ ), .ZN(\mexu/_0086_ ) );
OAI21_X1 \mexu/_1414_ ( .A(\mexu/_0990_ ), .B1(\mexu/_0595_ ), .B2(\mexu/_0596_ ), .ZN(\mexu/_0620_ ) );
BUF_X4 \mexu/_1415_ ( .A(\mexu/_0384_ ), .Z(\mexu/_0621_ ) );
NAND4_X1 \mexu/_1416_ ( .A1(\mexu/_0618_ ), .A2(\mexu/_1032_ ), .A3(\mexu/_0598_ ), .A4(\mexu/_0621_ ), .ZN(\mexu/_0622_ ) );
NAND2_X1 \mexu/_1417_ ( .A1(\mexu/_0620_ ), .A2(\mexu/_0622_ ), .ZN(\mexu/_0088_ ) );
BUF_X4 \mexu/_1418_ ( .A(\mexu/_0568_ ), .Z(\mexu/_0623_ ) );
BUF_X4 \mexu/_1419_ ( .A(\mexu/_0394_ ), .Z(\mexu/_0624_ ) );
OAI21_X1 \mexu/_1420_ ( .A(\mexu/_0991_ ), .B1(\mexu/_0623_ ), .B2(\mexu/_0624_ ), .ZN(\mexu/_0625_ ) );
BUF_X4 \mexu/_1421_ ( .A(\mexu/_0395_ ), .Z(\mexu/_0626_ ) );
NAND4_X1 \mexu/_1422_ ( .A1(\mexu/_0618_ ), .A2(\mexu/_1033_ ), .A3(\mexu/_0626_ ), .A4(\mexu/_0621_ ), .ZN(\mexu/_0627_ ) );
NAND2_X1 \mexu/_1423_ ( .A1(\mexu/_0625_ ), .A2(\mexu/_0627_ ), .ZN(\mexu/_0089_ ) );
OAI21_X1 \mexu/_1424_ ( .A(\mexu/_0992_ ), .B1(\mexu/_0623_ ), .B2(\mexu/_0624_ ), .ZN(\mexu/_0628_ ) );
NAND4_X1 \mexu/_1425_ ( .A1(\mexu/_0618_ ), .A2(\mexu/_1034_ ), .A3(\mexu/_0626_ ), .A4(\mexu/_0621_ ), .ZN(\mexu/_0629_ ) );
NAND2_X1 \mexu/_1426_ ( .A1(\mexu/_0628_ ), .A2(\mexu/_0629_ ), .ZN(\mexu/_0090_ ) );
OAI21_X1 \mexu/_1427_ ( .A(\mexu/_0993_ ), .B1(\mexu/_0623_ ), .B2(\mexu/_0624_ ), .ZN(\mexu/_0630_ ) );
NAND4_X1 \mexu/_1428_ ( .A1(\mexu/_0618_ ), .A2(\mexu/_1035_ ), .A3(\mexu/_0626_ ), .A4(\mexu/_0621_ ), .ZN(\mexu/_0631_ ) );
NAND2_X1 \mexu/_1429_ ( .A1(\mexu/_0630_ ), .A2(\mexu/_0631_ ), .ZN(\mexu/_0091_ ) );
OAI21_X1 \mexu/_1430_ ( .A(\mexu/_0994_ ), .B1(\mexu/_0623_ ), .B2(\mexu/_0624_ ), .ZN(\mexu/_0632_ ) );
NAND4_X1 \mexu/_1431_ ( .A1(\mexu/_0618_ ), .A2(\mexu/_1036_ ), .A3(\mexu/_0626_ ), .A4(\mexu/_0621_ ), .ZN(\mexu/_0633_ ) );
NAND2_X1 \mexu/_1432_ ( .A1(\mexu/_0632_ ), .A2(\mexu/_0633_ ), .ZN(\mexu/_0092_ ) );
OAI21_X1 \mexu/_1433_ ( .A(\mexu/_0995_ ), .B1(\mexu/_0623_ ), .B2(\mexu/_0624_ ), .ZN(\mexu/_0634_ ) );
NAND4_X1 \mexu/_1434_ ( .A1(\mexu/_0618_ ), .A2(\mexu/_1037_ ), .A3(\mexu/_0626_ ), .A4(\mexu/_0621_ ), .ZN(\mexu/_0635_ ) );
NAND2_X1 \mexu/_1435_ ( .A1(\mexu/_0634_ ), .A2(\mexu/_0635_ ), .ZN(\mexu/_0093_ ) );
OAI21_X1 \mexu/_1436_ ( .A(\mexu/_0996_ ), .B1(\mexu/_0623_ ), .B2(\mexu/_0624_ ), .ZN(\mexu/_0636_ ) );
NAND4_X1 \mexu/_1437_ ( .A1(\mexu/_0618_ ), .A2(\mexu/_1038_ ), .A3(\mexu/_0626_ ), .A4(\mexu/_0621_ ), .ZN(\mexu/_0637_ ) );
NAND2_X1 \mexu/_1438_ ( .A1(\mexu/_0636_ ), .A2(\mexu/_0637_ ), .ZN(\mexu/_0094_ ) );
OAI21_X1 \mexu/_1439_ ( .A(\mexu/_0997_ ), .B1(\mexu/_0623_ ), .B2(\mexu/_0624_ ), .ZN(\mexu/_0638_ ) );
NAND4_X1 \mexu/_1440_ ( .A1(\mexu/_0618_ ), .A2(\mexu/_1039_ ), .A3(\mexu/_0626_ ), .A4(\mexu/_0621_ ), .ZN(\mexu/_0639_ ) );
NAND2_X1 \mexu/_1441_ ( .A1(\mexu/_0638_ ), .A2(\mexu/_0639_ ), .ZN(\mexu/_0095_ ) );
OAI21_X1 \mexu/_1442_ ( .A(\mexu/_0998_ ), .B1(\mexu/_0623_ ), .B2(\mexu/_0624_ ), .ZN(\mexu/_0640_ ) );
NAND4_X1 \mexu/_1443_ ( .A1(\mexu/_0618_ ), .A2(\mexu/_1040_ ), .A3(\mexu/_0626_ ), .A4(\mexu/_0621_ ), .ZN(\mexu/_0641_ ) );
NAND2_X1 \mexu/_1444_ ( .A1(\mexu/_0640_ ), .A2(\mexu/_0641_ ), .ZN(\mexu/_0096_ ) );
OAI21_X1 \mexu/_1445_ ( .A(\mexu/_0999_ ), .B1(\mexu/_0623_ ), .B2(\mexu/_0624_ ), .ZN(\mexu/_0642_ ) );
NAND4_X1 \mexu/_1446_ ( .A1(\mexu/_0391_ ), .A2(\mexu/_1041_ ), .A3(\mexu/_0626_ ), .A4(\mexu/_0621_ ), .ZN(\mexu/_0643_ ) );
NAND2_X1 \mexu/_1447_ ( .A1(\mexu/_0642_ ), .A2(\mexu/_0643_ ), .ZN(\mexu/_0097_ ) );
OAI21_X1 \mexu/_1448_ ( .A(\mexu/_1001_ ), .B1(\mexu/_0623_ ), .B2(\mexu/_0624_ ), .ZN(\mexu/_0644_ ) );
NAND4_X1 \mexu/_1449_ ( .A1(\mexu/_0391_ ), .A2(\mexu/_1043_ ), .A3(\mexu/_0626_ ), .A4(\mexu/_0384_ ), .ZN(\mexu/_0645_ ) );
NAND2_X1 \mexu/_1450_ ( .A1(\mexu/_0644_ ), .A2(\mexu/_0645_ ), .ZN(\mexu/_0099_ ) );
OAI21_X1 \mexu/_1451_ ( .A(\mexu/_1002_ ), .B1(\mexu/_0568_ ), .B2(\mexu/_0394_ ), .ZN(\mexu/_0646_ ) );
NAND4_X1 \mexu/_1452_ ( .A1(\mexu/_0391_ ), .A2(\mexu/_1044_ ), .A3(\mexu/_0395_ ), .A4(\mexu/_0384_ ), .ZN(\mexu/_0647_ ) );
NAND2_X1 \mexu/_1453_ ( .A1(\mexu/_0646_ ), .A2(\mexu/_0647_ ), .ZN(\mexu/_0100_ ) );
NAND4_X1 \mexu/_1454_ ( .A1(\mexu/_0462_ ), .A2(\mexu/_0367_ ), .A3(\mexu/_0366_ ), .A4(\mexu/_0383_ ), .ZN(\mexu/_0648_ ) );
OAI21_X1 \mexu/_1455_ ( .A(\mexu/_0648_ ), .B1(\mexu/_0426_ ), .B2(\mexu/_0174_ ), .ZN(\mexu/_1019_ ) );
INV_X1 \mexu/_1456_ ( .A(\mexu/_0400_ ), .ZN(\mexu/_0649_ ) );
NOR4_X1 \mexu/_1457_ ( .A1(\mexu/_0175_ ), .A2(\mexu/_0173_ ), .A3(\mexu/_0174_ ), .A4(\mexu/_0203_ ), .ZN(\mexu/_0650_ ) );
NOR4_X1 \mexu/_1458_ ( .A1(\mexu/_0649_ ), .A2(\mexu/_0175_ ), .A3(\mexu/_0405_ ), .A4(\mexu/_0650_ ), .ZN(\mexu/_0651_ ) );
AND3_X1 \mexu/_1459_ ( .A1(\mexu/_0368_ ), .A2(\mexu/_0392_ ), .A3(\mexu/_0409_ ), .ZN(\mexu/_0652_ ) );
OR3_X1 \mexu/_1460_ ( .A1(\mexu/_0651_ ), .A2(\mexu/_0403_ ), .A3(\mexu/_0652_ ), .ZN(\mexu/_1084_ ) );
AND2_X1 \mexu/_1461_ ( .A1(\mexu/_0373_ ), .A2(\mexu/_0374_ ), .ZN(\mexu/_1018_ ) );
OAI21_X1 \mexu/_1462_ ( .A(\mexu/_0454_ ), .B1(\mexu/_0397_ ), .B2(\mexu/_0434_ ), .ZN(\mexu/_0208_ ) );
AND2_X4 \mexu/_1463_ ( .A1(\mexu/_0176_ ), .A2(\mexu/_0978_ ), .ZN(\mexu/_0653_ ) );
NOR2_X1 \mexu/_1464_ ( .A1(\mexu/_0176_ ), .A2(\mexu/_0978_ ), .ZN(\mexu/_0654_ ) );
AOI211_X4 \mexu/_1465_ ( .A(\mexu/_0653_ ), .B(\mexu/_0654_ ), .C1(\mexu/_0381_ ), .C2(\mexu/_0387_ ), .ZN(\mexu/_0039_ ) );
XOR2_X2 \mexu/_1466_ ( .A(\mexu/_0187_ ), .B(\mexu/_0989_ ), .Z(\mexu/_0655_ ) );
XOR2_X1 \mexu/_1467_ ( .A(\mexu/_0655_ ), .B(\mexu/_0653_ ), .Z(\mexu/_0656_ ) );
XOR2_X2 \mexu/_1468_ ( .A(\mexu/_0187_ ), .B(\mexu/_1031_ ), .Z(\mexu/_0657_ ) );
AND2_X4 \mexu/_1469_ ( .A1(\mexu/_0176_ ), .A2(\mexu/_1020_ ), .ZN(\mexu/_0658_ ) );
XOR2_X1 \mexu/_1470_ ( .A(\mexu/_0657_ ), .B(\mexu/_0658_ ), .Z(\mexu/_0659_ ) );
BUF_X4 \mexu/_1471_ ( .A(\mexu/_0388_ ), .Z(\mexu/_0660_ ) );
BUF_X4 \mexu/_1472_ ( .A(\mexu/_0660_ ), .Z(\mexu/_0661_ ) );
MUX2_X1 \mexu/_1473_ ( .A(\mexu/_0656_ ), .B(\mexu/_0659_ ), .S(\mexu/_0661_ ), .Z(\mexu/_0050_ ) );
AND2_X4 \mexu/_1474_ ( .A1(\mexu/_0655_ ), .A2(\mexu/_0653_ ), .ZN(\mexu/_0662_ ) );
AND2_X1 \mexu/_1475_ ( .A1(\mexu/_0187_ ), .A2(\mexu/_0989_ ), .ZN(\mexu/_0663_ ) );
NOR2_X4 \mexu/_1476_ ( .A1(\mexu/_0662_ ), .A2(\mexu/_0663_ ), .ZN(\mexu/_0664_ ) );
XOR2_X1 \mexu/_1477_ ( .A(\mexu/_0198_ ), .B(\mexu/_1000_ ), .Z(\mexu/_0665_ ) );
INV_X1 \mexu/_1478_ ( .A(\mexu/_0665_ ), .ZN(\mexu/_0666_ ) );
XNOR2_X1 \mexu/_1479_ ( .A(\mexu/_0664_ ), .B(\mexu/_0666_ ), .ZN(\mexu/_0667_ ) );
BUF_X4 \mexu/_1480_ ( .A(\mexu/_0661_ ), .Z(\mexu/_0668_ ) );
AND2_X4 \mexu/_1481_ ( .A1(\mexu/_0657_ ), .A2(\mexu/_0658_ ), .ZN(\mexu/_0669_ ) );
AND2_X1 \mexu/_1482_ ( .A1(\mexu/_0187_ ), .A2(\mexu/_1031_ ), .ZN(\mexu/_0670_ ) );
NOR2_X1 \mexu/_1483_ ( .A1(\mexu/_0669_ ), .A2(\mexu/_0670_ ), .ZN(\mexu/_0671_ ) );
INV_X1 \mexu/_1484_ ( .A(\mexu/_0671_ ), .ZN(\mexu/_0672_ ) );
XOR2_X2 \mexu/_1485_ ( .A(\mexu/_0198_ ), .B(\mexu/_1042_ ), .Z(\mexu/_0673_ ) );
AND2_X1 \mexu/_1486_ ( .A1(\mexu/_0672_ ), .A2(\mexu/_0673_ ), .ZN(\mexu/_0674_ ) );
OAI21_X1 \mexu/_1487_ ( .A(\mexu/_0661_ ), .B1(\mexu/_0672_ ), .B2(\mexu/_0673_ ), .ZN(\mexu/_0675_ ) );
OAI22_X1 \mexu/_1488_ ( .A1(\mexu/_0667_ ), .A2(\mexu/_0668_ ), .B1(\mexu/_0674_ ), .B2(\mexu/_0675_ ), .ZN(\mexu/_0061_ ) );
NOR2_X1 \mexu/_1489_ ( .A1(\mexu/_0664_ ), .A2(\mexu/_0666_ ), .ZN(\mexu/_0676_ ) );
AND2_X1 \mexu/_1490_ ( .A1(\mexu/_0198_ ), .A2(\mexu/_1000_ ), .ZN(\mexu/_0677_ ) );
NOR2_X1 \mexu/_1491_ ( .A1(\mexu/_0676_ ), .A2(\mexu/_0677_ ), .ZN(\mexu/_0678_ ) );
XOR2_X2 \mexu/_1492_ ( .A(\mexu/_0201_ ), .B(\mexu/_1003_ ), .Z(\mexu/_0679_ ) );
XNOR2_X1 \mexu/_1493_ ( .A(\mexu/_0678_ ), .B(\mexu/_0679_ ), .ZN(\mexu/_0680_ ) );
AND2_X1 \mexu/_1494_ ( .A1(\mexu/_0198_ ), .A2(\mexu/_1042_ ), .ZN(\mexu/_0681_ ) );
NOR2_X1 \mexu/_1495_ ( .A1(\mexu/_0674_ ), .A2(\mexu/_0681_ ), .ZN(\mexu/_0682_ ) );
XOR2_X2 \mexu/_1496_ ( .A(\mexu/_0201_ ), .B(\mexu/_1045_ ), .Z(\mexu/_0683_ ) );
XNOR2_X1 \mexu/_1497_ ( .A(\mexu/_0682_ ), .B(\mexu/_0683_ ), .ZN(\mexu/_0684_ ) );
MUX2_X1 \mexu/_1498_ ( .A(\mexu/_0680_ ), .B(\mexu/_0684_ ), .S(\mexu/_0661_ ), .Z(\mexu/_0064_ ) );
AND2_X2 \mexu/_1499_ ( .A1(\mexu/_0679_ ), .A2(\mexu/_0677_ ), .ZN(\mexu/_0685_ ) );
AOI21_X4 \mexu/_1500_ ( .A(\mexu/_0685_ ), .B1(\mexu/_0201_ ), .B2(\mexu/_1003_ ), .ZN(\mexu/_0686_ ) );
INV_X2 \mexu/_1501_ ( .A(\mexu/_0686_ ), .ZN(\mexu/_0687_ ) );
NAND2_X1 \mexu/_1502_ ( .A1(\mexu/_0665_ ), .A2(\mexu/_0679_ ), .ZN(\mexu/_0688_ ) );
NOR2_X4 \mexu/_1503_ ( .A1(\mexu/_0664_ ), .A2(\mexu/_0688_ ), .ZN(\mexu/_0689_ ) );
NOR2_X1 \mexu/_1504_ ( .A1(\mexu/_0687_ ), .A2(\mexu/_0689_ ), .ZN(\mexu/_0690_ ) );
XOR2_X2 \mexu/_1505_ ( .A(\mexu/_0202_ ), .B(\mexu/_1004_ ), .Z(\mexu/_0691_ ) );
INV_X1 \mexu/_1506_ ( .A(\mexu/_0691_ ), .ZN(\mexu/_0692_ ) );
XNOR2_X1 \mexu/_1507_ ( .A(\mexu/_0690_ ), .B(\mexu/_0692_ ), .ZN(\mexu/_0693_ ) );
AND2_X2 \mexu/_1508_ ( .A1(\mexu/_0683_ ), .A2(\mexu/_0681_ ), .ZN(\mexu/_0694_ ) );
AOI21_X4 \mexu/_1509_ ( .A(\mexu/_0694_ ), .B1(\mexu/_0201_ ), .B2(\mexu/_1045_ ), .ZN(\mexu/_0695_ ) );
OAI211_X2 \mexu/_1510_ ( .A(\mexu/_0673_ ), .B(\mexu/_0683_ ), .C1(\mexu/_0669_ ), .C2(\mexu/_0670_ ), .ZN(\mexu/_0696_ ) );
AND2_X4 \mexu/_1511_ ( .A1(\mexu/_0695_ ), .A2(\mexu/_0696_ ), .ZN(\mexu/_0697_ ) );
INV_X4 \mexu/_1512_ ( .A(\mexu/_0697_ ), .ZN(\mexu/_0698_ ) );
XOR2_X1 \mexu/_1513_ ( .A(\mexu/_0202_ ), .B(\mexu/_1046_ ), .Z(\mexu/_0699_ ) );
AND2_X1 \mexu/_1514_ ( .A1(\mexu/_0698_ ), .A2(\mexu/_0699_ ), .ZN(\mexu/_0700_ ) );
OAI21_X1 \mexu/_1515_ ( .A(\mexu/_0661_ ), .B1(\mexu/_0698_ ), .B2(\mexu/_0699_ ), .ZN(\mexu/_0701_ ) );
OAI22_X1 \mexu/_1516_ ( .A1(\mexu/_0693_ ), .A2(\mexu/_0668_ ), .B1(\mexu/_0700_ ), .B2(\mexu/_0701_ ), .ZN(\mexu/_0065_ ) );
NOR2_X1 \mexu/_1517_ ( .A1(\mexu/_0690_ ), .A2(\mexu/_0692_ ), .ZN(\mexu/_0702_ ) );
AND2_X1 \mexu/_1518_ ( .A1(\mexu/_0202_ ), .A2(\mexu/_1004_ ), .ZN(\mexu/_0703_ ) );
NOR2_X1 \mexu/_1519_ ( .A1(\mexu/_0702_ ), .A2(\mexu/_0703_ ), .ZN(\mexu/_0704_ ) );
AND2_X4 \mexu/_1520_ ( .A1(\mexu/_0203_ ), .A2(\mexu/_1005_ ), .ZN(\mexu/_0705_ ) );
NOR2_X4 \mexu/_1521_ ( .A1(\mexu/_0203_ ), .A2(\mexu/_1005_ ), .ZN(\mexu/_0706_ ) );
NOR2_X4 \mexu/_1522_ ( .A1(\mexu/_0705_ ), .A2(\mexu/_0706_ ), .ZN(\mexu/_0707_ ) );
XNOR2_X1 \mexu/_1523_ ( .A(\mexu/_0704_ ), .B(\mexu/_0707_ ), .ZN(\mexu/_0708_ ) );
AND2_X1 \mexu/_1524_ ( .A1(\mexu/_0202_ ), .A2(\mexu/_1046_ ), .ZN(\mexu/_0709_ ) );
NOR2_X1 \mexu/_1525_ ( .A1(\mexu/_0700_ ), .A2(\mexu/_0709_ ), .ZN(\mexu/_0710_ ) );
XOR2_X2 \mexu/_1526_ ( .A(\mexu/_0203_ ), .B(\mexu/_1047_ ), .Z(\mexu/_0711_ ) );
XNOR2_X1 \mexu/_1527_ ( .A(\mexu/_0710_ ), .B(\mexu/_0711_ ), .ZN(\mexu/_0712_ ) );
MUX2_X1 \mexu/_1528_ ( .A(\mexu/_0708_ ), .B(\mexu/_0712_ ), .S(\mexu/_0661_ ), .Z(\mexu/_0066_ ) );
XOR2_X2 \mexu/_1529_ ( .A(\mexu/_0204_ ), .B(\mexu/_1048_ ), .Z(\mexu/_0713_ ) );
INV_X1 \mexu/_1530_ ( .A(\mexu/_0713_ ), .ZN(\mexu/_0714_ ) );
AND2_X1 \mexu/_1531_ ( .A1(\mexu/_0699_ ), .A2(\mexu/_0711_ ), .ZN(\mexu/_0715_ ) );
NAND2_X1 \mexu/_1532_ ( .A1(\mexu/_0698_ ), .A2(\mexu/_0715_ ), .ZN(\mexu/_0716_ ) );
AND2_X4 \mexu/_1533_ ( .A1(\mexu/_0711_ ), .A2(\mexu/_0709_ ), .ZN(\mexu/_0717_ ) );
AOI21_X4 \mexu/_1534_ ( .A(\mexu/_0717_ ), .B1(\mexu/_0203_ ), .B2(\mexu/_1047_ ), .ZN(\mexu/_0718_ ) );
AOI21_X1 \mexu/_1535_ ( .A(\mexu/_0714_ ), .B1(\mexu/_0716_ ), .B2(\mexu/_0718_ ), .ZN(\mexu/_0719_ ) );
INV_X1 \mexu/_1536_ ( .A(\mexu/_0719_ ), .ZN(\mexu/_0720_ ) );
BUF_X4 \mexu/_1537_ ( .A(\mexu/_0660_ ), .Z(\mexu/_0721_ ) );
NAND3_X1 \mexu/_1538_ ( .A1(\mexu/_0716_ ), .A2(\mexu/_0714_ ), .A3(\mexu/_0718_ ), .ZN(\mexu/_0722_ ) );
NAND3_X1 \mexu/_1539_ ( .A1(\mexu/_0720_ ), .A2(\mexu/_0721_ ), .A3(\mexu/_0722_ ), .ZN(\mexu/_0723_ ) );
OAI211_X2 \mexu/_1540_ ( .A(\mexu/_0691_ ), .B(\mexu/_0707_ ), .C1(\mexu/_0687_ ), .C2(\mexu/_0689_ ), .ZN(\mexu/_0724_ ) );
AOI21_X2 \mexu/_1541_ ( .A(\mexu/_0705_ ), .B1(\mexu/_0707_ ), .B2(\mexu/_0703_ ), .ZN(\mexu/_0725_ ) );
XOR2_X2 \mexu/_1542_ ( .A(\mexu/_0204_ ), .B(\mexu/_1006_ ), .Z(\mexu/_0726_ ) );
INV_X1 \mexu/_1543_ ( .A(\mexu/_0726_ ), .ZN(\mexu/_0727_ ) );
AND3_X1 \mexu/_1544_ ( .A1(\mexu/_0724_ ), .A2(\mexu/_0725_ ), .A3(\mexu/_0727_ ), .ZN(\mexu/_0728_ ) );
AOI21_X1 \mexu/_1545_ ( .A(\mexu/_0727_ ), .B1(\mexu/_0724_ ), .B2(\mexu/_0725_ ), .ZN(\mexu/_0729_ ) );
OR3_X1 \mexu/_1546_ ( .A1(\mexu/_0728_ ), .A2(\mexu/_0729_ ), .A3(\mexu/_0660_ ), .ZN(\mexu/_0730_ ) );
NAND2_X1 \mexu/_1547_ ( .A1(\mexu/_0723_ ), .A2(\mexu/_0730_ ), .ZN(\mexu/_0067_ ) );
AND2_X1 \mexu/_1548_ ( .A1(\mexu/_0204_ ), .A2(\mexu/_1006_ ), .ZN(\mexu/_0731_ ) );
NOR2_X1 \mexu/_1549_ ( .A1(\mexu/_0729_ ), .A2(\mexu/_0731_ ), .ZN(\mexu/_0732_ ) );
XOR2_X2 \mexu/_1550_ ( .A(\mexu/_0205_ ), .B(\mexu/_1007_ ), .Z(\mexu/_0733_ ) );
INV_X1 \mexu/_1551_ ( .A(\mexu/_0733_ ), .ZN(\mexu/_0734_ ) );
XNOR2_X1 \mexu/_1552_ ( .A(\mexu/_0732_ ), .B(\mexu/_0734_ ), .ZN(\mexu/_0735_ ) );
NAND2_X1 \mexu/_1553_ ( .A1(\mexu/_0204_ ), .A2(\mexu/_1048_ ), .ZN(\mexu/_0736_ ) );
AND2_X4 \mexu/_1554_ ( .A1(\mexu/_0205_ ), .A2(\mexu/_1049_ ), .ZN(\mexu/_0737_ ) );
NOR2_X1 \mexu/_1555_ ( .A1(\mexu/_0205_ ), .A2(\mexu/_1049_ ), .ZN(\mexu/_0738_ ) );
NOR2_X2 \mexu/_1556_ ( .A1(\mexu/_0737_ ), .A2(\mexu/_0738_ ), .ZN(\mexu/_0739_ ) );
INV_X1 \mexu/_1557_ ( .A(\mexu/_0739_ ), .ZN(\mexu/_0740_ ) );
NAND3_X1 \mexu/_1558_ ( .A1(\mexu/_0720_ ), .A2(\mexu/_0736_ ), .A3(\mexu/_0740_ ), .ZN(\mexu/_0741_ ) );
BUF_X4 \mexu/_1559_ ( .A(\mexu/_0660_ ), .Z(\mexu/_0742_ ) );
NAND2_X1 \mexu/_1560_ ( .A1(\mexu/_0741_ ), .A2(\mexu/_0742_ ), .ZN(\mexu/_0743_ ) );
AOI21_X1 \mexu/_1561_ ( .A(\mexu/_0740_ ), .B1(\mexu/_0720_ ), .B2(\mexu/_0736_ ), .ZN(\mexu/_0744_ ) );
OAI22_X1 \mexu/_1562_ ( .A1(\mexu/_0735_ ), .A2(\mexu/_0668_ ), .B1(\mexu/_0743_ ), .B2(\mexu/_0744_ ), .ZN(\mexu/_0068_ ) );
NAND4_X4 \mexu/_1563_ ( .A1(\mexu/_0698_ ), .A2(\mexu/_0713_ ), .A3(\mexu/_0715_ ), .A4(\mexu/_0739_ ), .ZN(\mexu/_0745_ ) );
NOR3_X1 \mexu/_1564_ ( .A1(\mexu/_0718_ ), .A2(\mexu/_0714_ ), .A3(\mexu/_0740_ ), .ZN(\mexu/_0746_ ) );
NOR3_X1 \mexu/_1565_ ( .A1(\mexu/_0737_ ), .A2(\mexu/_0738_ ), .A3(\mexu/_0736_ ), .ZN(\mexu/_0747_ ) );
NOR3_X2 \mexu/_1566_ ( .A1(\mexu/_0746_ ), .A2(\mexu/_0737_ ), .A3(\mexu/_0747_ ), .ZN(\mexu/_0748_ ) );
AND2_X4 \mexu/_1567_ ( .A1(\mexu/_0745_ ), .A2(\mexu/_0748_ ), .ZN(\mexu/_0749_ ) );
INV_X4 \mexu/_1568_ ( .A(\mexu/_0749_ ), .ZN(\mexu/_0750_ ) );
XOR2_X1 \mexu/_1569_ ( .A(\mexu/_0206_ ), .B(\mexu/_1050_ ), .Z(\mexu/_0751_ ) );
OAI21_X1 \mexu/_1570_ ( .A(\mexu/_0721_ ), .B1(\mexu/_0750_ ), .B2(\mexu/_0751_ ), .ZN(\mexu/_0752_ ) );
AND2_X1 \mexu/_1571_ ( .A1(\mexu/_0206_ ), .A2(\mexu/_1050_ ), .ZN(\mexu/_0753_ ) );
NOR2_X1 \mexu/_1572_ ( .A1(\mexu/_0206_ ), .A2(\mexu/_1050_ ), .ZN(\mexu/_0754_ ) );
NOR3_X1 \mexu/_1573_ ( .A1(\mexu/_0749_ ), .A2(\mexu/_0753_ ), .A3(\mexu/_0754_ ), .ZN(\mexu/_0755_ ) );
AND2_X1 \mexu/_1574_ ( .A1(\mexu/_0733_ ), .A2(\mexu/_0731_ ), .ZN(\mexu/_0756_ ) );
NOR3_X2 \mexu/_1575_ ( .A1(\mexu/_0725_ ), .A2(\mexu/_0727_ ), .A3(\mexu/_0734_ ), .ZN(\mexu/_0757_ ) );
AOI211_X2 \mexu/_1576_ ( .A(\mexu/_0756_ ), .B(\mexu/_0757_ ), .C1(\mexu/_0205_ ), .C2(\mexu/_1007_ ), .ZN(\mexu/_0758_ ) );
AND4_X1 \mexu/_1577_ ( .A1(\mexu/_0691_ ), .A2(\mexu/_0726_ ), .A3(\mexu/_0733_ ), .A4(\mexu/_0707_ ), .ZN(\mexu/_0759_ ) );
OAI21_X2 \mexu/_1578_ ( .A(\mexu/_0759_ ), .B1(\mexu/_0687_ ), .B2(\mexu/_0689_ ), .ZN(\mexu/_0760_ ) );
AND2_X4 \mexu/_1579_ ( .A1(\mexu/_0758_ ), .A2(\mexu/_0760_ ), .ZN(\mexu/_0761_ ) );
XOR2_X1 \mexu/_1580_ ( .A(\mexu/_0206_ ), .B(\mexu/_1008_ ), .Z(\mexu/_0762_ ) );
INV_X1 \mexu/_1581_ ( .A(\mexu/_0762_ ), .ZN(\mexu/_0763_ ) );
XNOR2_X1 \mexu/_1582_ ( .A(\mexu/_0761_ ), .B(\mexu/_0763_ ), .ZN(\mexu/_0764_ ) );
OAI22_X1 \mexu/_1583_ ( .A1(\mexu/_0752_ ), .A2(\mexu/_0755_ ), .B1(\mexu/_0668_ ), .B2(\mexu/_0764_ ), .ZN(\mexu/_0069_ ) );
OR2_X1 \mexu/_1584_ ( .A1(\mexu/_0755_ ), .A2(\mexu/_0753_ ), .ZN(\mexu/_0765_ ) );
XOR2_X2 \mexu/_1585_ ( .A(\mexu/_0207_ ), .B(\mexu/_1051_ ), .Z(\mexu/_0766_ ) );
AND2_X1 \mexu/_1586_ ( .A1(\mexu/_0765_ ), .A2(\mexu/_0766_ ), .ZN(\mexu/_0767_ ) );
OAI21_X1 \mexu/_1587_ ( .A(\mexu/_0742_ ), .B1(\mexu/_0765_ ), .B2(\mexu/_0766_ ), .ZN(\mexu/_0768_ ) );
AOI21_X1 \mexu/_1588_ ( .A(\mexu/_0763_ ), .B1(\mexu/_0758_ ), .B2(\mexu/_0760_ ), .ZN(\mexu/_0769_ ) );
AND2_X1 \mexu/_1589_ ( .A1(\mexu/_0206_ ), .A2(\mexu/_1008_ ), .ZN(\mexu/_0770_ ) );
NOR2_X1 \mexu/_1590_ ( .A1(\mexu/_0769_ ), .A2(\mexu/_0770_ ), .ZN(\mexu/_0771_ ) );
AND2_X4 \mexu/_1591_ ( .A1(\mexu/_0207_ ), .A2(\mexu/_1009_ ), .ZN(\mexu/_0772_ ) );
NOR2_X1 \mexu/_1592_ ( .A1(\mexu/_0207_ ), .A2(\mexu/_1009_ ), .ZN(\mexu/_0773_ ) );
NOR2_X2 \mexu/_1593_ ( .A1(\mexu/_0772_ ), .A2(\mexu/_0773_ ), .ZN(\mexu/_0774_ ) );
XOR2_X1 \mexu/_1594_ ( .A(\mexu/_0771_ ), .B(\mexu/_0774_ ), .Z(\mexu/_0775_ ) );
BUF_X4 \mexu/_1595_ ( .A(\mexu/_0661_ ), .Z(\mexu/_0776_ ) );
OAI22_X1 \mexu/_1596_ ( .A1(\mexu/_0767_ ), .A2(\mexu/_0768_ ), .B1(\mexu/_0775_ ), .B2(\mexu/_0776_ ), .ZN(\mexu/_0070_ ) );
INV_X4 \mexu/_1597_ ( .A(\mexu/_0761_ ), .ZN(\mexu/_0777_ ) );
AND2_X1 \mexu/_1598_ ( .A1(\mexu/_0762_ ), .A2(\mexu/_0774_ ), .ZN(\mexu/_0778_ ) );
NAND2_X1 \mexu/_1599_ ( .A1(\mexu/_0777_ ), .A2(\mexu/_0778_ ), .ZN(\mexu/_0779_ ) );
AOI21_X1 \mexu/_1600_ ( .A(\mexu/_0772_ ), .B1(\mexu/_0774_ ), .B2(\mexu/_0770_ ), .ZN(\mexu/_0780_ ) );
XOR2_X1 \mexu/_1601_ ( .A(\mexu/_0177_ ), .B(\mexu/_0979_ ), .Z(\mexu/_0781_ ) );
INV_X1 \mexu/_1602_ ( .A(\mexu/_0781_ ), .ZN(\mexu/_0782_ ) );
AND3_X1 \mexu/_1603_ ( .A1(\mexu/_0779_ ), .A2(\mexu/_0780_ ), .A3(\mexu/_0782_ ), .ZN(\mexu/_0783_ ) );
AOI21_X1 \mexu/_1604_ ( .A(\mexu/_0782_ ), .B1(\mexu/_0779_ ), .B2(\mexu/_0780_ ), .ZN(\mexu/_0784_ ) );
OR3_X1 \mexu/_1605_ ( .A1(\mexu/_0783_ ), .A2(\mexu/_0784_ ), .A3(\mexu/_0660_ ), .ZN(\mexu/_0785_ ) );
AND2_X1 \mexu/_1606_ ( .A1(\mexu/_0751_ ), .A2(\mexu/_0766_ ), .ZN(\mexu/_0786_ ) );
NAND2_X1 \mexu/_1607_ ( .A1(\mexu/_0750_ ), .A2(\mexu/_0786_ ), .ZN(\mexu/_0787_ ) );
AND2_X2 \mexu/_1608_ ( .A1(\mexu/_0766_ ), .A2(\mexu/_0753_ ), .ZN(\mexu/_0788_ ) );
AOI21_X2 \mexu/_1609_ ( .A(\mexu/_0788_ ), .B1(\mexu/_0207_ ), .B2(\mexu/_1051_ ), .ZN(\mexu/_0789_ ) );
AND2_X1 \mexu/_1610_ ( .A1(\mexu/_0787_ ), .A2(\mexu/_0789_ ), .ZN(\mexu/_0790_ ) );
XOR2_X1 \mexu/_1611_ ( .A(\mexu/_0177_ ), .B(\mexu/_1021_ ), .Z(\mexu/_0791_ ) );
INV_X1 \mexu/_1612_ ( .A(\mexu/_0791_ ), .ZN(\mexu/_0792_ ) );
XNOR2_X1 \mexu/_1613_ ( .A(\mexu/_0790_ ), .B(\mexu/_0792_ ), .ZN(\mexu/_0793_ ) );
INV_X1 \mexu/_1614_ ( .A(\mexu/_0660_ ), .ZN(\mexu/_0794_ ) );
OAI21_X1 \mexu/_1615_ ( .A(\mexu/_0785_ ), .B1(\mexu/_0793_ ), .B2(\mexu/_0794_ ), .ZN(\mexu/_0040_ ) );
XOR2_X1 \mexu/_1616_ ( .A(\mexu/_0178_ ), .B(\mexu/_1022_ ), .Z(\mexu/_0795_ ) );
INV_X1 \mexu/_1617_ ( .A(\mexu/_0795_ ), .ZN(\mexu/_0796_ ) );
OR2_X1 \mexu/_1618_ ( .A1(\mexu/_0790_ ), .A2(\mexu/_0792_ ), .ZN(\mexu/_0797_ ) );
NAND2_X1 \mexu/_1619_ ( .A1(\mexu/_0177_ ), .A2(\mexu/_1021_ ), .ZN(\mexu/_0798_ ) );
AOI21_X1 \mexu/_1620_ ( .A(\mexu/_0796_ ), .B1(\mexu/_0797_ ), .B2(\mexu/_0798_ ), .ZN(\mexu/_0799_ ) );
OAI211_X2 \mexu/_1621_ ( .A(\mexu/_0798_ ), .B(\mexu/_0796_ ), .C1(\mexu/_0790_ ), .C2(\mexu/_0792_ ), .ZN(\mexu/_0800_ ) );
NAND2_X1 \mexu/_1622_ ( .A1(\mexu/_0800_ ), .A2(\mexu/_0721_ ), .ZN(\mexu/_0801_ ) );
AND2_X1 \mexu/_1623_ ( .A1(\mexu/_0177_ ), .A2(\mexu/_0979_ ), .ZN(\mexu/_0802_ ) );
NOR2_X1 \mexu/_1624_ ( .A1(\mexu/_0784_ ), .A2(\mexu/_0802_ ), .ZN(\mexu/_0803_ ) );
XOR2_X1 \mexu/_1625_ ( .A(\mexu/_0178_ ), .B(\mexu/_0980_ ), .Z(\mexu/_0804_ ) );
INV_X1 \mexu/_1626_ ( .A(\mexu/_0804_ ), .ZN(\mexu/_0805_ ) );
XNOR2_X1 \mexu/_1627_ ( .A(\mexu/_0803_ ), .B(\mexu/_0805_ ), .ZN(\mexu/_0806_ ) );
OAI22_X1 \mexu/_1628_ ( .A1(\mexu/_0799_ ), .A2(\mexu/_0801_ ), .B1(\mexu/_0668_ ), .B2(\mexu/_0806_ ), .ZN(\mexu/_0041_ ) );
XOR2_X1 \mexu/_1629_ ( .A(\mexu/_0179_ ), .B(\mexu/_1023_ ), .Z(\mexu/_0807_ ) );
INV_X1 \mexu/_1630_ ( .A(\mexu/_0807_ ), .ZN(\mexu/_0808_ ) );
AND3_X1 \mexu/_1631_ ( .A1(\mexu/_0786_ ), .A2(\mexu/_0791_ ), .A3(\mexu/_0795_ ), .ZN(\mexu/_0809_ ) );
NAND2_X1 \mexu/_1632_ ( .A1(\mexu/_0750_ ), .A2(\mexu/_0809_ ), .ZN(\mexu/_0810_ ) );
NOR3_X2 \mexu/_1633_ ( .A1(\mexu/_0789_ ), .A2(\mexu/_0792_ ), .A3(\mexu/_0796_ ), .ZN(\mexu/_0811_ ) );
AND2_X1 \mexu/_1634_ ( .A1(\mexu/_0178_ ), .A2(\mexu/_1022_ ), .ZN(\mexu/_0812_ ) );
AND3_X1 \mexu/_1635_ ( .A1(\mexu/_0795_ ), .A2(\mexu/_0177_ ), .A3(\mexu/_1021_ ), .ZN(\mexu/_0813_ ) );
NOR3_X4 \mexu/_1636_ ( .A1(\mexu/_0811_ ), .A2(\mexu/_0812_ ), .A3(\mexu/_0813_ ), .ZN(\mexu/_0814_ ) );
AOI21_X1 \mexu/_1637_ ( .A(\mexu/_0808_ ), .B1(\mexu/_0810_ ), .B2(\mexu/_0814_ ), .ZN(\mexu/_0815_ ) );
INV_X1 \mexu/_1638_ ( .A(\mexu/_0815_ ), .ZN(\mexu/_0816_ ) );
NAND3_X1 \mexu/_1639_ ( .A1(\mexu/_0810_ ), .A2(\mexu/_0814_ ), .A3(\mexu/_0808_ ), .ZN(\mexu/_0817_ ) );
NAND3_X1 \mexu/_1640_ ( .A1(\mexu/_0816_ ), .A2(\mexu/_0721_ ), .A3(\mexu/_0817_ ), .ZN(\mexu/_0818_ ) );
AND3_X1 \mexu/_1641_ ( .A1(\mexu/_0778_ ), .A2(\mexu/_0781_ ), .A3(\mexu/_0804_ ), .ZN(\mexu/_0819_ ) );
NAND2_X1 \mexu/_1642_ ( .A1(\mexu/_0777_ ), .A2(\mexu/_0819_ ), .ZN(\mexu/_0820_ ) );
NOR3_X2 \mexu/_1643_ ( .A1(\mexu/_0780_ ), .A2(\mexu/_0782_ ), .A3(\mexu/_0805_ ), .ZN(\mexu/_0821_ ) );
AND2_X1 \mexu/_1644_ ( .A1(\mexu/_0178_ ), .A2(\mexu/_0980_ ), .ZN(\mexu/_0822_ ) );
AND2_X1 \mexu/_1645_ ( .A1(\mexu/_0804_ ), .A2(\mexu/_0802_ ), .ZN(\mexu/_0823_ ) );
NOR3_X2 \mexu/_1646_ ( .A1(\mexu/_0821_ ), .A2(\mexu/_0822_ ), .A3(\mexu/_0823_ ), .ZN(\mexu/_0824_ ) );
AND2_X1 \mexu/_1647_ ( .A1(\mexu/_0820_ ), .A2(\mexu/_0824_ ), .ZN(\mexu/_0825_ ) );
XOR2_X1 \mexu/_1648_ ( .A(\mexu/_0179_ ), .B(\mexu/_0981_ ), .Z(\mexu/_0826_ ) );
INV_X1 \mexu/_1649_ ( .A(\mexu/_0826_ ), .ZN(\mexu/_0827_ ) );
XNOR2_X1 \mexu/_1650_ ( .A(\mexu/_0825_ ), .B(\mexu/_0827_ ), .ZN(\mexu/_0828_ ) );
OAI21_X1 \mexu/_1651_ ( .A(\mexu/_0818_ ), .B1(\mexu/_0828_ ), .B2(\mexu/_0668_ ), .ZN(\mexu/_0042_ ) );
AOI21_X1 \mexu/_1652_ ( .A(\mexu/_0827_ ), .B1(\mexu/_0820_ ), .B2(\mexu/_0824_ ), .ZN(\mexu/_0829_ ) );
AND2_X1 \mexu/_1653_ ( .A1(\mexu/_0179_ ), .A2(\mexu/_0981_ ), .ZN(\mexu/_0830_ ) );
NOR2_X1 \mexu/_1654_ ( .A1(\mexu/_0829_ ), .A2(\mexu/_0830_ ), .ZN(\mexu/_0831_ ) );
AND2_X4 \mexu/_1655_ ( .A1(\mexu/_0180_ ), .A2(\mexu/_0982_ ), .ZN(\mexu/_0832_ ) );
NOR2_X1 \mexu/_1656_ ( .A1(\mexu/_0180_ ), .A2(\mexu/_0982_ ), .ZN(\mexu/_0833_ ) );
NOR2_X2 \mexu/_1657_ ( .A1(\mexu/_0832_ ), .A2(\mexu/_0833_ ), .ZN(\mexu/_0834_ ) );
XNOR2_X1 \mexu/_1658_ ( .A(\mexu/_0831_ ), .B(\mexu/_0834_ ), .ZN(\mexu/_0835_ ) );
AND2_X1 \mexu/_1659_ ( .A1(\mexu/_0179_ ), .A2(\mexu/_1023_ ), .ZN(\mexu/_0836_ ) );
NOR2_X1 \mexu/_1660_ ( .A1(\mexu/_0815_ ), .A2(\mexu/_0836_ ), .ZN(\mexu/_0837_ ) );
AND2_X4 \mexu/_1661_ ( .A1(\mexu/_0180_ ), .A2(\mexu/_1024_ ), .ZN(\mexu/_0838_ ) );
NOR2_X1 \mexu/_1662_ ( .A1(\mexu/_0180_ ), .A2(\mexu/_1024_ ), .ZN(\mexu/_0839_ ) );
NOR2_X1 \mexu/_1663_ ( .A1(\mexu/_0838_ ), .A2(\mexu/_0839_ ), .ZN(\mexu/_0840_ ) );
XNOR2_X1 \mexu/_1664_ ( .A(\mexu/_0837_ ), .B(\mexu/_0840_ ), .ZN(\mexu/_0841_ ) );
MUX2_X1 \mexu/_1665_ ( .A(\mexu/_0835_ ), .B(\mexu/_0841_ ), .S(\mexu/_0661_ ), .Z(\mexu/_0043_ ) );
INV_X1 \mexu/_1666_ ( .A(\mexu/_0836_ ), .ZN(\mexu/_0842_ ) );
AOI21_X1 \mexu/_1667_ ( .A(\mexu/_0839_ ), .B1(\mexu/_0816_ ), .B2(\mexu/_0842_ ), .ZN(\mexu/_0843_ ) );
XOR2_X1 \mexu/_1668_ ( .A(\mexu/_0181_ ), .B(\mexu/_1025_ ), .Z(\mexu/_0844_ ) );
OR3_X1 \mexu/_1669_ ( .A1(\mexu/_0843_ ), .A2(\mexu/_0838_ ), .A3(\mexu/_0844_ ), .ZN(\mexu/_0845_ ) );
OAI21_X1 \mexu/_1670_ ( .A(\mexu/_0844_ ), .B1(\mexu/_0843_ ), .B2(\mexu/_0838_ ), .ZN(\mexu/_0846_ ) );
NAND3_X1 \mexu/_1671_ ( .A1(\mexu/_0845_ ), .A2(\mexu/_0721_ ), .A3(\mexu/_0846_ ), .ZN(\mexu/_0847_ ) );
AND2_X2 \mexu/_1672_ ( .A1(\mexu/_0826_ ), .A2(\mexu/_0834_ ), .ZN(\mexu/_0848_ ) );
INV_X1 \mexu/_1673_ ( .A(\mexu/_0848_ ), .ZN(\mexu/_0849_ ) );
OR2_X1 \mexu/_1674_ ( .A1(\mexu/_0825_ ), .A2(\mexu/_0849_ ), .ZN(\mexu/_0850_ ) );
XOR2_X1 \mexu/_1675_ ( .A(\mexu/_0181_ ), .B(\mexu/_0983_ ), .Z(\mexu/_0851_ ) );
INV_X1 \mexu/_1676_ ( .A(\mexu/_0851_ ), .ZN(\mexu/_0852_ ) );
AOI21_X1 \mexu/_1677_ ( .A(\mexu/_0832_ ), .B1(\mexu/_0834_ ), .B2(\mexu/_0830_ ), .ZN(\mexu/_0853_ ) );
AND3_X1 \mexu/_1678_ ( .A1(\mexu/_0850_ ), .A2(\mexu/_0852_ ), .A3(\mexu/_0853_ ), .ZN(\mexu/_0854_ ) );
AOI21_X1 \mexu/_1679_ ( .A(\mexu/_0852_ ), .B1(\mexu/_0850_ ), .B2(\mexu/_0853_ ), .ZN(\mexu/_0855_ ) );
OR3_X1 \mexu/_1680_ ( .A1(\mexu/_0854_ ), .A2(\mexu/_0855_ ), .A3(\mexu/_0660_ ), .ZN(\mexu/_0856_ ) );
NAND2_X1 \mexu/_1681_ ( .A1(\mexu/_0847_ ), .A2(\mexu/_0856_ ), .ZN(\mexu/_0044_ ) );
NAND2_X1 \mexu/_1682_ ( .A1(\mexu/_0181_ ), .A2(\mexu/_1025_ ), .ZN(\mexu/_0857_ ) );
NAND2_X1 \mexu/_1683_ ( .A1(\mexu/_0846_ ), .A2(\mexu/_0857_ ), .ZN(\mexu/_0858_ ) );
XOR2_X2 \mexu/_1684_ ( .A(\mexu/_0182_ ), .B(\mexu/_1026_ ), .Z(\mexu/_0859_ ) );
AND2_X1 \mexu/_1685_ ( .A1(\mexu/_0858_ ), .A2(\mexu/_0859_ ), .ZN(\mexu/_0860_ ) );
OAI21_X1 \mexu/_1686_ ( .A(\mexu/_0742_ ), .B1(\mexu/_0858_ ), .B2(\mexu/_0859_ ), .ZN(\mexu/_0861_ ) );
AND2_X1 \mexu/_1687_ ( .A1(\mexu/_0181_ ), .A2(\mexu/_0983_ ), .ZN(\mexu/_0862_ ) );
NOR2_X1 \mexu/_1688_ ( .A1(\mexu/_0855_ ), .A2(\mexu/_0862_ ), .ZN(\mexu/_0863_ ) );
XOR2_X2 \mexu/_1689_ ( .A(\mexu/_0182_ ), .B(\mexu/_0984_ ), .Z(\mexu/_0864_ ) );
INV_X1 \mexu/_1690_ ( .A(\mexu/_0864_ ), .ZN(\mexu/_0865_ ) );
XNOR2_X1 \mexu/_1691_ ( .A(\mexu/_0863_ ), .B(\mexu/_0865_ ), .ZN(\mexu/_0866_ ) );
OAI22_X1 \mexu/_1692_ ( .A1(\mexu/_0860_ ), .A2(\mexu/_0861_ ), .B1(\mexu/_0866_ ), .B2(\mexu/_0776_ ), .ZN(\mexu/_0045_ ) );
AND2_X2 \mexu/_1693_ ( .A1(\mexu/_0844_ ), .A2(\mexu/_0859_ ), .ZN(\mexu/_0867_ ) );
AND2_X1 \mexu/_1694_ ( .A1(\mexu/_0807_ ), .A2(\mexu/_0840_ ), .ZN(\mexu/_0868_ ) );
AND2_X1 \mexu/_1695_ ( .A1(\mexu/_0867_ ), .A2(\mexu/_0868_ ), .ZN(\mexu/_0869_ ) );
NAND3_X2 \mexu/_1696_ ( .A1(\mexu/_0750_ ), .A2(\mexu/_0809_ ), .A3(\mexu/_0869_ ), .ZN(\mexu/_0870_ ) );
NAND3_X1 \mexu/_1697_ ( .A1(\mexu/_0859_ ), .A2(\mexu/_0181_ ), .A3(\mexu/_1025_ ), .ZN(\mexu/_0871_ ) );
INV_X1 \mexu/_1698_ ( .A(\mexu/_0869_ ), .ZN(\mexu/_0872_ ) );
OAI221_X1 \mexu/_1699_ ( .A(\mexu/_0871_ ), .B1(\mexu/_0509_ ), .B2(\mexu/_0610_ ), .C1(\mexu/_0814_ ), .C2(\mexu/_0872_ ), .ZN(\mexu/_0873_ ) );
INV_X1 \mexu/_1700_ ( .A(\mexu/_0838_ ), .ZN(\mexu/_0874_ ) );
AOI21_X1 \mexu/_1701_ ( .A(\mexu/_0839_ ), .B1(\mexu/_0842_ ), .B2(\mexu/_0874_ ), .ZN(\mexu/_0875_ ) );
AOI21_X1 \mexu/_1702_ ( .A(\mexu/_0873_ ), .B1(\mexu/_0875_ ), .B2(\mexu/_0867_ ), .ZN(\mexu/_0876_ ) );
AND2_X2 \mexu/_1703_ ( .A1(\mexu/_0870_ ), .A2(\mexu/_0876_ ), .ZN(\mexu/_0877_ ) );
INV_X4 \mexu/_1704_ ( .A(\mexu/_0877_ ), .ZN(\mexu/_0878_ ) );
XOR2_X1 \mexu/_1705_ ( .A(\mexu/_0183_ ), .B(\mexu/_1027_ ), .Z(\mexu/_0879_ ) );
OAI21_X1 \mexu/_1706_ ( .A(\mexu/_0742_ ), .B1(\mexu/_0878_ ), .B2(\mexu/_0879_ ), .ZN(\mexu/_0880_ ) );
AND2_X1 \mexu/_1707_ ( .A1(\mexu/_0183_ ), .A2(\mexu/_1027_ ), .ZN(\mexu/_0881_ ) );
NOR2_X1 \mexu/_1708_ ( .A1(\mexu/_0183_ ), .A2(\mexu/_1027_ ), .ZN(\mexu/_0882_ ) );
NOR3_X1 \mexu/_1709_ ( .A1(\mexu/_0877_ ), .A2(\mexu/_0881_ ), .A3(\mexu/_0882_ ), .ZN(\mexu/_0883_ ) );
AND2_X1 \mexu/_1710_ ( .A1(\mexu/_0851_ ), .A2(\mexu/_0864_ ), .ZN(\mexu/_0884_ ) );
AND2_X2 \mexu/_1711_ ( .A1(\mexu/_0884_ ), .A2(\mexu/_0848_ ), .ZN(\mexu/_0885_ ) );
NAND3_X4 \mexu/_1712_ ( .A1(\mexu/_0777_ ), .A2(\mexu/_0819_ ), .A3(\mexu/_0885_ ), .ZN(\mexu/_0886_ ) );
INV_X1 \mexu/_1713_ ( .A(\mexu/_0885_ ), .ZN(\mexu/_0887_ ) );
NOR2_X2 \mexu/_1714_ ( .A1(\mexu/_0824_ ), .A2(\mexu/_0887_ ), .ZN(\mexu/_0888_ ) );
AND2_X1 \mexu/_1715_ ( .A1(\mexu/_0182_ ), .A2(\mexu/_0984_ ), .ZN(\mexu/_0889_ ) );
NOR3_X1 \mexu/_1716_ ( .A1(\mexu/_0853_ ), .A2(\mexu/_0852_ ), .A3(\mexu/_0865_ ), .ZN(\mexu/_0890_ ) );
AND2_X1 \mexu/_1717_ ( .A1(\mexu/_0864_ ), .A2(\mexu/_0862_ ), .ZN(\mexu/_0891_ ) );
NOR4_X4 \mexu/_1718_ ( .A1(\mexu/_0888_ ), .A2(\mexu/_0889_ ), .A3(\mexu/_0890_ ), .A4(\mexu/_0891_ ), .ZN(\mexu/_0892_ ) );
AND2_X4 \mexu/_1719_ ( .A1(\mexu/_0886_ ), .A2(\mexu/_0892_ ), .ZN(\mexu/_0893_ ) );
XOR2_X1 \mexu/_1720_ ( .A(\mexu/_0183_ ), .B(\mexu/_0985_ ), .Z(\mexu/_0894_ ) );
INV_X1 \mexu/_1721_ ( .A(\mexu/_0894_ ), .ZN(\mexu/_0895_ ) );
XNOR2_X1 \mexu/_1722_ ( .A(\mexu/_0893_ ), .B(\mexu/_0895_ ), .ZN(\mexu/_0896_ ) );
OAI22_X1 \mexu/_1723_ ( .A1(\mexu/_0880_ ), .A2(\mexu/_0883_ ), .B1(\mexu/_0668_ ), .B2(\mexu/_0896_ ), .ZN(\mexu/_0046_ ) );
OR2_X1 \mexu/_1724_ ( .A1(\mexu/_0883_ ), .A2(\mexu/_0881_ ), .ZN(\mexu/_0897_ ) );
XOR2_X1 \mexu/_1725_ ( .A(\mexu/_0184_ ), .B(\mexu/_1028_ ), .Z(\mexu/_0898_ ) );
AND2_X1 \mexu/_1726_ ( .A1(\mexu/_0897_ ), .A2(\mexu/_0898_ ), .ZN(\mexu/_0899_ ) );
OAI21_X1 \mexu/_1727_ ( .A(\mexu/_0742_ ), .B1(\mexu/_0897_ ), .B2(\mexu/_0898_ ), .ZN(\mexu/_0900_ ) );
AOI21_X1 \mexu/_1728_ ( .A(\mexu/_0895_ ), .B1(\mexu/_0886_ ), .B2(\mexu/_0892_ ), .ZN(\mexu/_0901_ ) );
AND2_X1 \mexu/_1729_ ( .A1(\mexu/_0183_ ), .A2(\mexu/_0985_ ), .ZN(\mexu/_0902_ ) );
NOR2_X1 \mexu/_1730_ ( .A1(\mexu/_0901_ ), .A2(\mexu/_0902_ ), .ZN(\mexu/_0903_ ) );
AND2_X1 \mexu/_1731_ ( .A1(\mexu/_0184_ ), .A2(\mexu/_0986_ ), .ZN(\mexu/_0904_ ) );
NOR2_X1 \mexu/_1732_ ( .A1(\mexu/_0184_ ), .A2(\mexu/_0986_ ), .ZN(\mexu/_0905_ ) );
NOR2_X1 \mexu/_1733_ ( .A1(\mexu/_0904_ ), .A2(\mexu/_0905_ ), .ZN(\mexu/_0906_ ) );
XOR2_X1 \mexu/_1734_ ( .A(\mexu/_0903_ ), .B(\mexu/_0906_ ), .Z(\mexu/_0907_ ) );
OAI22_X1 \mexu/_1735_ ( .A1(\mexu/_0899_ ), .A2(\mexu/_0900_ ), .B1(\mexu/_0776_ ), .B2(\mexu/_0907_ ), .ZN(\mexu/_0047_ ) );
INV_X4 \mexu/_1736_ ( .A(\mexu/_0893_ ), .ZN(\mexu/_0908_ ) );
AND2_X1 \mexu/_1737_ ( .A1(\mexu/_0894_ ), .A2(\mexu/_0906_ ), .ZN(\mexu/_0909_ ) );
NAND2_X1 \mexu/_1738_ ( .A1(\mexu/_0908_ ), .A2(\mexu/_0909_ ), .ZN(\mexu/_0910_ ) );
AOI21_X1 \mexu/_1739_ ( .A(\mexu/_0904_ ), .B1(\mexu/_0906_ ), .B2(\mexu/_0902_ ), .ZN(\mexu/_0911_ ) );
XOR2_X1 \mexu/_1740_ ( .A(\mexu/_0185_ ), .B(\mexu/_0987_ ), .Z(\mexu/_0912_ ) );
INV_X1 \mexu/_1741_ ( .A(\mexu/_0912_ ), .ZN(\mexu/_0913_ ) );
AND3_X1 \mexu/_1742_ ( .A1(\mexu/_0910_ ), .A2(\mexu/_0911_ ), .A3(\mexu/_0913_ ), .ZN(\mexu/_0914_ ) );
AOI21_X1 \mexu/_1743_ ( .A(\mexu/_0913_ ), .B1(\mexu/_0910_ ), .B2(\mexu/_0911_ ), .ZN(\mexu/_0915_ ) );
OR3_X1 \mexu/_1744_ ( .A1(\mexu/_0914_ ), .A2(\mexu/_0915_ ), .A3(\mexu/_0660_ ), .ZN(\mexu/_0916_ ) );
AND2_X1 \mexu/_1745_ ( .A1(\mexu/_0879_ ), .A2(\mexu/_0898_ ), .ZN(\mexu/_0917_ ) );
NAND2_X1 \mexu/_1746_ ( .A1(\mexu/_0878_ ), .A2(\mexu/_0917_ ), .ZN(\mexu/_0918_ ) );
AND2_X1 \mexu/_1747_ ( .A1(\mexu/_0898_ ), .A2(\mexu/_0881_ ), .ZN(\mexu/_0919_ ) );
AOI21_X1 \mexu/_1748_ ( .A(\mexu/_0919_ ), .B1(\mexu/_0184_ ), .B2(\mexu/_1028_ ), .ZN(\mexu/_0920_ ) );
AND2_X1 \mexu/_1749_ ( .A1(\mexu/_0918_ ), .A2(\mexu/_0920_ ), .ZN(\mexu/_0921_ ) );
XOR2_X1 \mexu/_1750_ ( .A(\mexu/_0185_ ), .B(\mexu/_1029_ ), .Z(\mexu/_0922_ ) );
INV_X1 \mexu/_1751_ ( .A(\mexu/_0922_ ), .ZN(\mexu/_0923_ ) );
XNOR2_X1 \mexu/_1752_ ( .A(\mexu/_0921_ ), .B(\mexu/_0923_ ), .ZN(\mexu/_0924_ ) );
OAI21_X1 \mexu/_1753_ ( .A(\mexu/_0916_ ), .B1(\mexu/_0924_ ), .B2(\mexu/_0794_ ), .ZN(\mexu/_0048_ ) );
XOR2_X1 \mexu/_1754_ ( .A(\mexu/_0186_ ), .B(\mexu/_1030_ ), .Z(\mexu/_0925_ ) );
INV_X1 \mexu/_1755_ ( .A(\mexu/_0925_ ), .ZN(\mexu/_0926_ ) );
OR2_X1 \mexu/_1756_ ( .A1(\mexu/_0921_ ), .A2(\mexu/_0923_ ), .ZN(\mexu/_0927_ ) );
NAND2_X1 \mexu/_1757_ ( .A1(\mexu/_0185_ ), .A2(\mexu/_1029_ ), .ZN(\mexu/_0928_ ) );
AOI21_X1 \mexu/_1758_ ( .A(\mexu/_0926_ ), .B1(\mexu/_0927_ ), .B2(\mexu/_0928_ ), .ZN(\mexu/_0929_ ) );
OAI211_X2 \mexu/_1759_ ( .A(\mexu/_0928_ ), .B(\mexu/_0926_ ), .C1(\mexu/_0921_ ), .C2(\mexu/_0923_ ), .ZN(\mexu/_0930_ ) );
NAND2_X1 \mexu/_1760_ ( .A1(\mexu/_0930_ ), .A2(\mexu/_0721_ ), .ZN(\mexu/_0931_ ) );
AND2_X1 \mexu/_1761_ ( .A1(\mexu/_0185_ ), .A2(\mexu/_0987_ ), .ZN(\mexu/_0932_ ) );
NOR2_X1 \mexu/_1762_ ( .A1(\mexu/_0915_ ), .A2(\mexu/_0932_ ), .ZN(\mexu/_0933_ ) );
XOR2_X1 \mexu/_1763_ ( .A(\mexu/_0186_ ), .B(\mexu/_0988_ ), .Z(\mexu/_0934_ ) );
INV_X1 \mexu/_1764_ ( .A(\mexu/_0934_ ), .ZN(\mexu/_0935_ ) );
XNOR2_X1 \mexu/_1765_ ( .A(\mexu/_0933_ ), .B(\mexu/_0935_ ), .ZN(\mexu/_0936_ ) );
OAI22_X1 \mexu/_1766_ ( .A1(\mexu/_0929_ ), .A2(\mexu/_0931_ ), .B1(\mexu/_0776_ ), .B2(\mexu/_0936_ ), .ZN(\mexu/_0049_ ) );
AND3_X1 \mexu/_1767_ ( .A1(\mexu/_0917_ ), .A2(\mexu/_0922_ ), .A3(\mexu/_0925_ ), .ZN(\mexu/_0937_ ) );
NAND2_X1 \mexu/_1768_ ( .A1(\mexu/_0878_ ), .A2(\mexu/_0937_ ), .ZN(\mexu/_0938_ ) );
NOR3_X1 \mexu/_1769_ ( .A1(\mexu/_0920_ ), .A2(\mexu/_0923_ ), .A3(\mexu/_0926_ ), .ZN(\mexu/_0939_ ) );
AND2_X1 \mexu/_1770_ ( .A1(\mexu/_0186_ ), .A2(\mexu/_1030_ ), .ZN(\mexu/_0940_ ) );
AND3_X1 \mexu/_1771_ ( .A1(\mexu/_0925_ ), .A2(\mexu/_0185_ ), .A3(\mexu/_1029_ ), .ZN(\mexu/_0941_ ) );
NOR3_X1 \mexu/_1772_ ( .A1(\mexu/_0939_ ), .A2(\mexu/_0940_ ), .A3(\mexu/_0941_ ), .ZN(\mexu/_0942_ ) );
AND2_X2 \mexu/_1773_ ( .A1(\mexu/_0938_ ), .A2(\mexu/_0942_ ), .ZN(\mexu/_0943_ ) );
INV_X1 \mexu/_1774_ ( .A(\mexu/_0943_ ), .ZN(\mexu/_0944_ ) );
XOR2_X1 \mexu/_1775_ ( .A(\mexu/_0188_ ), .B(\mexu/_1032_ ), .Z(\mexu/_0945_ ) );
AND2_X1 \mexu/_1776_ ( .A1(\mexu/_0944_ ), .A2(\mexu/_0945_ ), .ZN(\mexu/_0946_ ) );
OAI21_X1 \mexu/_1777_ ( .A(\mexu/_0742_ ), .B1(\mexu/_0944_ ), .B2(\mexu/_0945_ ), .ZN(\mexu/_0947_ ) );
AND3_X1 \mexu/_1778_ ( .A1(\mexu/_0909_ ), .A2(\mexu/_0912_ ), .A3(\mexu/_0934_ ), .ZN(\mexu/_0948_ ) );
NAND2_X1 \mexu/_1779_ ( .A1(\mexu/_0908_ ), .A2(\mexu/_0948_ ), .ZN(\mexu/_0949_ ) );
NOR3_X1 \mexu/_1780_ ( .A1(\mexu/_0911_ ), .A2(\mexu/_0913_ ), .A3(\mexu/_0935_ ), .ZN(\mexu/_0950_ ) );
AND2_X1 \mexu/_1781_ ( .A1(\mexu/_0186_ ), .A2(\mexu/_0988_ ), .ZN(\mexu/_0951_ ) );
AND2_X1 \mexu/_1782_ ( .A1(\mexu/_0934_ ), .A2(\mexu/_0932_ ), .ZN(\mexu/_0952_ ) );
NOR3_X1 \mexu/_1783_ ( .A1(\mexu/_0950_ ), .A2(\mexu/_0951_ ), .A3(\mexu/_0952_ ), .ZN(\mexu/_0953_ ) );
AND2_X1 \mexu/_1784_ ( .A1(\mexu/_0949_ ), .A2(\mexu/_0953_ ), .ZN(\mexu/_0954_ ) );
XOR2_X1 \mexu/_1785_ ( .A(\mexu/_0188_ ), .B(\mexu/_0990_ ), .Z(\mexu/_0955_ ) );
INV_X1 \mexu/_1786_ ( .A(\mexu/_0955_ ), .ZN(\mexu/_0956_ ) );
XNOR2_X1 \mexu/_1787_ ( .A(\mexu/_0954_ ), .B(\mexu/_0956_ ), .ZN(\mexu/_0957_ ) );
OAI22_X1 \mexu/_1788_ ( .A1(\mexu/_0946_ ), .A2(\mexu/_0947_ ), .B1(\mexu/_0776_ ), .B2(\mexu/_0957_ ), .ZN(\mexu/_0051_ ) );
AND2_X1 \mexu/_1789_ ( .A1(\mexu/_0188_ ), .A2(\mexu/_1032_ ), .ZN(\mexu/_0958_ ) );
XOR2_X1 \mexu/_1790_ ( .A(\mexu/_0189_ ), .B(\mexu/_1033_ ), .Z(\mexu/_0959_ ) );
OR3_X1 \mexu/_1791_ ( .A1(\mexu/_0946_ ), .A2(\mexu/_0958_ ), .A3(\mexu/_0959_ ), .ZN(\mexu/_0960_ ) );
OAI21_X1 \mexu/_1792_ ( .A(\mexu/_0959_ ), .B1(\mexu/_0946_ ), .B2(\mexu/_0958_ ), .ZN(\mexu/_0961_ ) );
NAND3_X1 \mexu/_1793_ ( .A1(\mexu/_0960_ ), .A2(\mexu/_0721_ ), .A3(\mexu/_0961_ ), .ZN(\mexu/_0962_ ) );
AOI21_X1 \mexu/_1794_ ( .A(\mexu/_0956_ ), .B1(\mexu/_0949_ ), .B2(\mexu/_0953_ ), .ZN(\mexu/_0963_ ) );
AND2_X1 \mexu/_1795_ ( .A1(\mexu/_0188_ ), .A2(\mexu/_0990_ ), .ZN(\mexu/_0964_ ) );
NOR2_X1 \mexu/_1796_ ( .A1(\mexu/_0963_ ), .A2(\mexu/_0964_ ), .ZN(\mexu/_0965_ ) );
XOR2_X2 \mexu/_1797_ ( .A(\mexu/_0189_ ), .B(\mexu/_0991_ ), .Z(\mexu/_0966_ ) );
XOR2_X1 \mexu/_1798_ ( .A(\mexu/_0965_ ), .B(\mexu/_0966_ ), .Z(\mexu/_0967_ ) );
OAI21_X1 \mexu/_1799_ ( .A(\mexu/_0962_ ), .B1(\mexu/_0668_ ), .B2(\mexu/_0967_ ), .ZN(\mexu/_0052_ ) );
AND2_X1 \mexu/_1800_ ( .A1(\mexu/_0955_ ), .A2(\mexu/_0966_ ), .ZN(\mexu/_0968_ ) );
INV_X1 \mexu/_1801_ ( .A(\mexu/_0968_ ), .ZN(\mexu/_0969_ ) );
OR2_X1 \mexu/_1802_ ( .A1(\mexu/_0954_ ), .A2(\mexu/_0969_ ), .ZN(\mexu/_0970_ ) );
XOR2_X1 \mexu/_1803_ ( .A(\mexu/_0190_ ), .B(\mexu/_0992_ ), .Z(\mexu/_0214_ ) );
INV_X1 \mexu/_1804_ ( .A(\mexu/_0214_ ), .ZN(\mexu/_0215_ ) );
AND2_X1 \mexu/_1805_ ( .A1(\mexu/_0966_ ), .A2(\mexu/_0964_ ), .ZN(\mexu/_0216_ ) );
AOI21_X1 \mexu/_1806_ ( .A(\mexu/_0216_ ), .B1(\mexu/_0189_ ), .B2(\mexu/_0991_ ), .ZN(\mexu/_0217_ ) );
AND3_X1 \mexu/_1807_ ( .A1(\mexu/_0970_ ), .A2(\mexu/_0215_ ), .A3(\mexu/_0217_ ), .ZN(\mexu/_0218_ ) );
AOI21_X1 \mexu/_1808_ ( .A(\mexu/_0215_ ), .B1(\mexu/_0970_ ), .B2(\mexu/_0217_ ), .ZN(\mexu/_0219_ ) );
OR3_X1 \mexu/_1809_ ( .A1(\mexu/_0218_ ), .A2(\mexu/_0219_ ), .A3(\mexu/_0660_ ), .ZN(\mexu/_0220_ ) );
AND2_X1 \mexu/_1810_ ( .A1(\mexu/_0945_ ), .A2(\mexu/_0959_ ), .ZN(\mexu/_0221_ ) );
INV_X1 \mexu/_1811_ ( .A(\mexu/_0221_ ), .ZN(\mexu/_0222_ ) );
OR2_X1 \mexu/_1812_ ( .A1(\mexu/_0943_ ), .A2(\mexu/_0222_ ), .ZN(\mexu/_0223_ ) );
AND2_X1 \mexu/_1813_ ( .A1(\mexu/_0959_ ), .A2(\mexu/_0958_ ), .ZN(\mexu/_0224_ ) );
AOI21_X1 \mexu/_1814_ ( .A(\mexu/_0224_ ), .B1(\mexu/_0189_ ), .B2(\mexu/_1033_ ), .ZN(\mexu/_0225_ ) );
NAND2_X1 \mexu/_1815_ ( .A1(\mexu/_0223_ ), .A2(\mexu/_0225_ ), .ZN(\mexu/_0226_ ) );
XOR2_X1 \mexu/_1816_ ( .A(\mexu/_0190_ ), .B(\mexu/_1034_ ), .Z(\mexu/_0227_ ) );
AND2_X2 \mexu/_1817_ ( .A1(\mexu/_0226_ ), .A2(\mexu/_0227_ ), .ZN(\mexu/_0228_ ) );
OAI21_X1 \mexu/_1818_ ( .A(\mexu/_0742_ ), .B1(\mexu/_0226_ ), .B2(\mexu/_0227_ ), .ZN(\mexu/_0229_ ) );
OAI21_X1 \mexu/_1819_ ( .A(\mexu/_0220_ ), .B1(\mexu/_0228_ ), .B2(\mexu/_0229_ ), .ZN(\mexu/_0053_ ) );
INV_X1 \mexu/_1820_ ( .A(\mexu/_0228_ ), .ZN(\mexu/_0230_ ) );
NAND2_X1 \mexu/_1821_ ( .A1(\mexu/_0190_ ), .A2(\mexu/_1034_ ), .ZN(\mexu/_0231_ ) );
AND2_X2 \mexu/_1822_ ( .A1(\mexu/_0191_ ), .A2(\mexu/_1035_ ), .ZN(\mexu/_0232_ ) );
NOR2_X1 \mexu/_1823_ ( .A1(\mexu/_0191_ ), .A2(\mexu/_1035_ ), .ZN(\mexu/_0233_ ) );
OAI211_X2 \mexu/_1824_ ( .A(\mexu/_0230_ ), .B(\mexu/_0231_ ), .C1(\mexu/_0232_ ), .C2(\mexu/_0233_ ), .ZN(\mexu/_0234_ ) );
NAND2_X1 \mexu/_1825_ ( .A1(\mexu/_0234_ ), .A2(\mexu/_0721_ ), .ZN(\mexu/_0235_ ) );
AOI211_X2 \mexu/_1826_ ( .A(\mexu/_0232_ ), .B(\mexu/_0233_ ), .C1(\mexu/_0230_ ), .C2(\mexu/_0231_ ), .ZN(\mexu/_0236_ ) );
AND2_X1 \mexu/_1827_ ( .A1(\mexu/_0190_ ), .A2(\mexu/_0992_ ), .ZN(\mexu/_0237_ ) );
NOR2_X1 \mexu/_1828_ ( .A1(\mexu/_0219_ ), .A2(\mexu/_0237_ ), .ZN(\mexu/_0238_ ) );
XOR2_X1 \mexu/_1829_ ( .A(\mexu/_0191_ ), .B(\mexu/_0993_ ), .Z(\mexu/_0239_ ) );
INV_X1 \mexu/_1830_ ( .A(\mexu/_0239_ ), .ZN(\mexu/_0240_ ) );
XNOR2_X1 \mexu/_1831_ ( .A(\mexu/_0238_ ), .B(\mexu/_0240_ ), .ZN(\mexu/_0241_ ) );
OAI22_X1 \mexu/_1832_ ( .A1(\mexu/_0235_ ), .A2(\mexu/_0236_ ), .B1(\mexu/_0241_ ), .B2(\mexu/_0776_ ), .ZN(\mexu/_0054_ ) );
NOR2_X1 \mexu/_1833_ ( .A1(\mexu/_0232_ ), .A2(\mexu/_0233_ ), .ZN(\mexu/_0242_ ) );
AND2_X1 \mexu/_1834_ ( .A1(\mexu/_0227_ ), .A2(\mexu/_0242_ ), .ZN(\mexu/_0243_ ) );
NAND4_X4 \mexu/_1835_ ( .A1(\mexu/_0878_ ), .A2(\mexu/_0937_ ), .A3(\mexu/_0221_ ), .A4(\mexu/_0243_ ), .ZN(\mexu/_0244_ ) );
INV_X1 \mexu/_1836_ ( .A(\mexu/_0243_ ), .ZN(\mexu/_0245_ ) );
NOR3_X1 \mexu/_1837_ ( .A1(\mexu/_0942_ ), .A2(\mexu/_0222_ ), .A3(\mexu/_0245_ ), .ZN(\mexu/_0246_ ) );
NOR2_X1 \mexu/_1838_ ( .A1(\mexu/_0225_ ), .A2(\mexu/_0245_ ), .ZN(\mexu/_0247_ ) );
NOR3_X1 \mexu/_1839_ ( .A1(\mexu/_0232_ ), .A2(\mexu/_0233_ ), .A3(\mexu/_0231_ ), .ZN(\mexu/_0248_ ) );
NOR4_X1 \mexu/_1840_ ( .A1(\mexu/_0246_ ), .A2(\mexu/_0232_ ), .A3(\mexu/_0247_ ), .A4(\mexu/_0248_ ), .ZN(\mexu/_0249_ ) );
AND2_X4 \mexu/_1841_ ( .A1(\mexu/_0244_ ), .A2(\mexu/_0249_ ), .ZN(\mexu/_0250_ ) );
INV_X4 \mexu/_1842_ ( .A(\mexu/_0250_ ), .ZN(\mexu/_0251_ ) );
XOR2_X1 \mexu/_1843_ ( .A(\mexu/_0192_ ), .B(\mexu/_1036_ ), .Z(\mexu/_0252_ ) );
OAI21_X1 \mexu/_1844_ ( .A(\mexu/_0742_ ), .B1(\mexu/_0251_ ), .B2(\mexu/_0252_ ), .ZN(\mexu/_0253_ ) );
AND2_X1 \mexu/_1845_ ( .A1(\mexu/_0192_ ), .A2(\mexu/_1036_ ), .ZN(\mexu/_0254_ ) );
NOR2_X1 \mexu/_1846_ ( .A1(\mexu/_0192_ ), .A2(\mexu/_1036_ ), .ZN(\mexu/_0255_ ) );
NOR3_X1 \mexu/_1847_ ( .A1(\mexu/_0250_ ), .A2(\mexu/_0254_ ), .A3(\mexu/_0255_ ), .ZN(\mexu/_0256_ ) );
AND2_X1 \mexu/_1848_ ( .A1(\mexu/_0214_ ), .A2(\mexu/_0239_ ), .ZN(\mexu/_0257_ ) );
NAND4_X4 \mexu/_1849_ ( .A1(\mexu/_0908_ ), .A2(\mexu/_0948_ ), .A3(\mexu/_0968_ ), .A4(\mexu/_0257_ ), .ZN(\mexu/_0258_ ) );
AND2_X1 \mexu/_1850_ ( .A1(\mexu/_0239_ ), .A2(\mexu/_0237_ ), .ZN(\mexu/_0259_ ) );
OR3_X2 \mexu/_1851_ ( .A1(\mexu/_0217_ ), .A2(\mexu/_0215_ ), .A3(\mexu/_0240_ ), .ZN(\mexu/_0260_ ) );
AND2_X1 \mexu/_1852_ ( .A1(\mexu/_0257_ ), .A2(\mexu/_0968_ ), .ZN(\mexu/_0261_ ) );
INV_X1 \mexu/_1853_ ( .A(\mexu/_0261_ ), .ZN(\mexu/_0262_ ) );
OAI21_X1 \mexu/_1854_ ( .A(\mexu/_0260_ ), .B1(\mexu/_0953_ ), .B2(\mexu/_0262_ ), .ZN(\mexu/_0263_ ) );
AOI211_X2 \mexu/_1855_ ( .A(\mexu/_0259_ ), .B(\mexu/_0263_ ), .C1(\mexu/_0191_ ), .C2(\mexu/_0993_ ), .ZN(\mexu/_0264_ ) );
AND2_X4 \mexu/_1856_ ( .A1(\mexu/_0258_ ), .A2(\mexu/_0264_ ), .ZN(\mexu/_0265_ ) );
XOR2_X1 \mexu/_1857_ ( .A(\mexu/_0192_ ), .B(\mexu/_0994_ ), .Z(\mexu/_0266_ ) );
INV_X1 \mexu/_1858_ ( .A(\mexu/_0266_ ), .ZN(\mexu/_0267_ ) );
XNOR2_X1 \mexu/_1859_ ( .A(\mexu/_0265_ ), .B(\mexu/_0267_ ), .ZN(\mexu/_0268_ ) );
OAI22_X1 \mexu/_1860_ ( .A1(\mexu/_0253_ ), .A2(\mexu/_0256_ ), .B1(\mexu/_0776_ ), .B2(\mexu/_0268_ ), .ZN(\mexu/_0055_ ) );
XOR2_X1 \mexu/_1861_ ( .A(\mexu/_0193_ ), .B(\mexu/_1037_ ), .Z(\mexu/_0269_ ) );
OR3_X1 \mexu/_1862_ ( .A1(\mexu/_0256_ ), .A2(\mexu/_0254_ ), .A3(\mexu/_0269_ ), .ZN(\mexu/_0270_ ) );
OAI21_X1 \mexu/_1863_ ( .A(\mexu/_0269_ ), .B1(\mexu/_0256_ ), .B2(\mexu/_0254_ ), .ZN(\mexu/_0271_ ) );
NAND3_X1 \mexu/_1864_ ( .A1(\mexu/_0270_ ), .A2(\mexu/_0721_ ), .A3(\mexu/_0271_ ), .ZN(\mexu/_0272_ ) );
AOI21_X1 \mexu/_1865_ ( .A(\mexu/_0267_ ), .B1(\mexu/_0258_ ), .B2(\mexu/_0264_ ), .ZN(\mexu/_0273_ ) );
AND2_X1 \mexu/_1866_ ( .A1(\mexu/_0192_ ), .A2(\mexu/_0994_ ), .ZN(\mexu/_0274_ ) );
NOR2_X1 \mexu/_1867_ ( .A1(\mexu/_0273_ ), .A2(\mexu/_0274_ ), .ZN(\mexu/_0275_ ) );
AND2_X1 \mexu/_1868_ ( .A1(\mexu/_0193_ ), .A2(\mexu/_0995_ ), .ZN(\mexu/_0276_ ) );
NOR2_X1 \mexu/_1869_ ( .A1(\mexu/_0193_ ), .A2(\mexu/_0995_ ), .ZN(\mexu/_0277_ ) );
NOR2_X1 \mexu/_1870_ ( .A1(\mexu/_0276_ ), .A2(\mexu/_0277_ ), .ZN(\mexu/_0278_ ) );
XOR2_X1 \mexu/_1871_ ( .A(\mexu/_0275_ ), .B(\mexu/_0278_ ), .Z(\mexu/_0279_ ) );
OAI21_X1 \mexu/_1872_ ( .A(\mexu/_0272_ ), .B1(\mexu/_0668_ ), .B2(\mexu/_0279_ ), .ZN(\mexu/_0056_ ) );
XOR2_X1 \mexu/_1873_ ( .A(\mexu/_0194_ ), .B(\mexu/_1038_ ), .Z(\mexu/_0280_ ) );
INV_X1 \mexu/_1874_ ( .A(\mexu/_0280_ ), .ZN(\mexu/_0281_ ) );
AND2_X1 \mexu/_1875_ ( .A1(\mexu/_0252_ ), .A2(\mexu/_0269_ ), .ZN(\mexu/_0282_ ) );
NAND2_X1 \mexu/_1876_ ( .A1(\mexu/_0251_ ), .A2(\mexu/_0282_ ), .ZN(\mexu/_0283_ ) );
AND2_X1 \mexu/_1877_ ( .A1(\mexu/_0269_ ), .A2(\mexu/_0254_ ), .ZN(\mexu/_0284_ ) );
AOI21_X1 \mexu/_1878_ ( .A(\mexu/_0284_ ), .B1(\mexu/_0193_ ), .B2(\mexu/_1037_ ), .ZN(\mexu/_0285_ ) );
AOI21_X1 \mexu/_1879_ ( .A(\mexu/_0281_ ), .B1(\mexu/_0283_ ), .B2(\mexu/_0285_ ), .ZN(\mexu/_0286_ ) );
INV_X1 \mexu/_1880_ ( .A(\mexu/_0286_ ), .ZN(\mexu/_0287_ ) );
NAND3_X1 \mexu/_1881_ ( .A1(\mexu/_0283_ ), .A2(\mexu/_0285_ ), .A3(\mexu/_0281_ ), .ZN(\mexu/_0288_ ) );
NAND3_X1 \mexu/_1882_ ( .A1(\mexu/_0287_ ), .A2(\mexu/_0721_ ), .A3(\mexu/_0288_ ), .ZN(\mexu/_0289_ ) );
XOR2_X1 \mexu/_1883_ ( .A(\mexu/_0194_ ), .B(\mexu/_0996_ ), .Z(\mexu/_0290_ ) );
INV_X1 \mexu/_1884_ ( .A(\mexu/_0290_ ), .ZN(\mexu/_0291_ ) );
INV_X4 \mexu/_1885_ ( .A(\mexu/_0265_ ), .ZN(\mexu/_0292_ ) );
AND2_X1 \mexu/_1886_ ( .A1(\mexu/_0266_ ), .A2(\mexu/_0278_ ), .ZN(\mexu/_0293_ ) );
NAND2_X1 \mexu/_1887_ ( .A1(\mexu/_0292_ ), .A2(\mexu/_0293_ ), .ZN(\mexu/_0294_ ) );
AOI21_X1 \mexu/_1888_ ( .A(\mexu/_0276_ ), .B1(\mexu/_0278_ ), .B2(\mexu/_0274_ ), .ZN(\mexu/_0295_ ) );
AOI21_X1 \mexu/_1889_ ( .A(\mexu/_0291_ ), .B1(\mexu/_0294_ ), .B2(\mexu/_0295_ ), .ZN(\mexu/_0296_ ) );
NAND3_X1 \mexu/_1890_ ( .A1(\mexu/_0294_ ), .A2(\mexu/_0291_ ), .A3(\mexu/_0295_ ), .ZN(\mexu/_0297_ ) );
NAND2_X1 \mexu/_1891_ ( .A1(\mexu/_0297_ ), .A2(\mexu/_0794_ ), .ZN(\mexu/_0298_ ) );
OAI21_X1 \mexu/_1892_ ( .A(\mexu/_0289_ ), .B1(\mexu/_0296_ ), .B2(\mexu/_0298_ ), .ZN(\mexu/_0057_ ) );
AND2_X1 \mexu/_1893_ ( .A1(\mexu/_0194_ ), .A2(\mexu/_0996_ ), .ZN(\mexu/_0299_ ) );
NOR2_X1 \mexu/_1894_ ( .A1(\mexu/_0296_ ), .A2(\mexu/_0299_ ), .ZN(\mexu/_0300_ ) );
XOR2_X1 \mexu/_1895_ ( .A(\mexu/_0195_ ), .B(\mexu/_0997_ ), .Z(\mexu/_0301_ ) );
INV_X1 \mexu/_1896_ ( .A(\mexu/_0301_ ), .ZN(\mexu/_0302_ ) );
XNOR2_X1 \mexu/_1897_ ( .A(\mexu/_0300_ ), .B(\mexu/_0302_ ), .ZN(\mexu/_0303_ ) );
XOR2_X1 \mexu/_1898_ ( .A(\mexu/_0195_ ), .B(\mexu/_1039_ ), .Z(\mexu/_0304_ ) );
AND2_X1 \mexu/_1899_ ( .A1(\mexu/_0194_ ), .A2(\mexu/_1038_ ), .ZN(\mexu/_0305_ ) );
OAI21_X1 \mexu/_1900_ ( .A(\mexu/_0304_ ), .B1(\mexu/_0286_ ), .B2(\mexu/_0305_ ), .ZN(\mexu/_0306_ ) );
NAND2_X1 \mexu/_1901_ ( .A1(\mexu/_0306_ ), .A2(\mexu/_0742_ ), .ZN(\mexu/_0307_ ) );
NOR3_X1 \mexu/_1902_ ( .A1(\mexu/_0286_ ), .A2(\mexu/_0305_ ), .A3(\mexu/_0304_ ), .ZN(\mexu/_0308_ ) );
OAI22_X1 \mexu/_1903_ ( .A1(\mexu/_0303_ ), .A2(\mexu/_0668_ ), .B1(\mexu/_0307_ ), .B2(\mexu/_0308_ ), .ZN(\mexu/_0058_ ) );
NAND4_X4 \mexu/_1904_ ( .A1(\mexu/_0251_ ), .A2(\mexu/_0282_ ), .A3(\mexu/_0280_ ), .A4(\mexu/_0304_ ), .ZN(\mexu/_0309_ ) );
AND2_X1 \mexu/_1905_ ( .A1(\mexu/_0304_ ), .A2(\mexu/_0305_ ), .ZN(\mexu/_0310_ ) );
INV_X1 \mexu/_1906_ ( .A(\mexu/_0285_ ), .ZN(\mexu/_0311_ ) );
AND3_X1 \mexu/_1907_ ( .A1(\mexu/_0311_ ), .A2(\mexu/_0280_ ), .A3(\mexu/_0304_ ), .ZN(\mexu/_0312_ ) );
AOI211_X4 \mexu/_1908_ ( .A(\mexu/_0310_ ), .B(\mexu/_0312_ ), .C1(\mexu/_0195_ ), .C2(\mexu/_1039_ ), .ZN(\mexu/_0313_ ) );
AND2_X4 \mexu/_1909_ ( .A1(\mexu/_0309_ ), .A2(\mexu/_0313_ ), .ZN(\mexu/_0314_ ) );
INV_X4 \mexu/_1910_ ( .A(\mexu/_0314_ ), .ZN(\mexu/_0315_ ) );
XOR2_X1 \mexu/_1911_ ( .A(\mexu/_0196_ ), .B(\mexu/_1040_ ), .Z(\mexu/_0316_ ) );
OAI21_X1 \mexu/_1912_ ( .A(\mexu/_0742_ ), .B1(\mexu/_0315_ ), .B2(\mexu/_0316_ ), .ZN(\mexu/_0317_ ) );
AND2_X1 \mexu/_1913_ ( .A1(\mexu/_0196_ ), .A2(\mexu/_1040_ ), .ZN(\mexu/_0318_ ) );
NOR2_X1 \mexu/_1914_ ( .A1(\mexu/_0196_ ), .A2(\mexu/_1040_ ), .ZN(\mexu/_0319_ ) );
NOR3_X1 \mexu/_1915_ ( .A1(\mexu/_0314_ ), .A2(\mexu/_0318_ ), .A3(\mexu/_0319_ ), .ZN(\mexu/_0320_ ) );
NAND4_X4 \mexu/_1916_ ( .A1(\mexu/_0292_ ), .A2(\mexu/_0290_ ), .A3(\mexu/_0293_ ), .A4(\mexu/_0301_ ), .ZN(\mexu/_0321_ ) );
AND2_X1 \mexu/_1917_ ( .A1(\mexu/_0301_ ), .A2(\mexu/_0299_ ), .ZN(\mexu/_0322_ ) );
NOR3_X1 \mexu/_1918_ ( .A1(\mexu/_0295_ ), .A2(\mexu/_0291_ ), .A3(\mexu/_0302_ ), .ZN(\mexu/_0323_ ) );
AOI211_X4 \mexu/_1919_ ( .A(\mexu/_0322_ ), .B(\mexu/_0323_ ), .C1(\mexu/_0195_ ), .C2(\mexu/_0997_ ), .ZN(\mexu/_0324_ ) );
AND2_X4 \mexu/_1920_ ( .A1(\mexu/_0321_ ), .A2(\mexu/_0324_ ), .ZN(\mexu/_0325_ ) );
XOR2_X1 \mexu/_1921_ ( .A(\mexu/_0196_ ), .B(\mexu/_0998_ ), .Z(\mexu/_0326_ ) );
INV_X1 \mexu/_1922_ ( .A(\mexu/_0326_ ), .ZN(\mexu/_0327_ ) );
XNOR2_X1 \mexu/_1923_ ( .A(\mexu/_0325_ ), .B(\mexu/_0327_ ), .ZN(\mexu/_0328_ ) );
OAI22_X1 \mexu/_1924_ ( .A1(\mexu/_0317_ ), .A2(\mexu/_0320_ ), .B1(\mexu/_0776_ ), .B2(\mexu/_0328_ ), .ZN(\mexu/_0059_ ) );
OR2_X1 \mexu/_1925_ ( .A1(\mexu/_0320_ ), .A2(\mexu/_0318_ ), .ZN(\mexu/_0329_ ) );
XOR2_X1 \mexu/_1926_ ( .A(\mexu/_0197_ ), .B(\mexu/_1041_ ), .Z(\mexu/_0330_ ) );
AND2_X1 \mexu/_1927_ ( .A1(\mexu/_0329_ ), .A2(\mexu/_0330_ ), .ZN(\mexu/_0331_ ) );
OAI21_X1 \mexu/_1928_ ( .A(\mexu/_0661_ ), .B1(\mexu/_0329_ ), .B2(\mexu/_0330_ ), .ZN(\mexu/_0332_ ) );
AOI21_X1 \mexu/_1929_ ( .A(\mexu/_0327_ ), .B1(\mexu/_0321_ ), .B2(\mexu/_0324_ ), .ZN(\mexu/_0333_ ) );
AND2_X1 \mexu/_1930_ ( .A1(\mexu/_0196_ ), .A2(\mexu/_0998_ ), .ZN(\mexu/_0334_ ) );
NOR2_X1 \mexu/_1931_ ( .A1(\mexu/_0333_ ), .A2(\mexu/_0334_ ), .ZN(\mexu/_0335_ ) );
AND2_X1 \mexu/_1932_ ( .A1(\mexu/_0197_ ), .A2(\mexu/_0999_ ), .ZN(\mexu/_0336_ ) );
NOR2_X1 \mexu/_1933_ ( .A1(\mexu/_0197_ ), .A2(\mexu/_0999_ ), .ZN(\mexu/_0337_ ) );
NOR2_X1 \mexu/_1934_ ( .A1(\mexu/_0336_ ), .A2(\mexu/_0337_ ), .ZN(\mexu/_0338_ ) );
XOR2_X1 \mexu/_1935_ ( .A(\mexu/_0335_ ), .B(\mexu/_0338_ ), .Z(\mexu/_0339_ ) );
OAI22_X1 \mexu/_1936_ ( .A1(\mexu/_0331_ ), .A2(\mexu/_0332_ ), .B1(\mexu/_0776_ ), .B2(\mexu/_0339_ ), .ZN(\mexu/_0060_ ) );
NAND3_X2 \mexu/_1937_ ( .A1(\mexu/_0315_ ), .A2(\mexu/_0316_ ), .A3(\mexu/_0330_ ), .ZN(\mexu/_0340_ ) );
AND2_X1 \mexu/_1938_ ( .A1(\mexu/_0330_ ), .A2(\mexu/_0318_ ), .ZN(\mexu/_0341_ ) );
AOI21_X1 \mexu/_1939_ ( .A(\mexu/_0341_ ), .B1(\mexu/_0197_ ), .B2(\mexu/_1041_ ), .ZN(\mexu/_0342_ ) );
AND2_X4 \mexu/_1940_ ( .A1(\mexu/_0340_ ), .A2(\mexu/_0342_ ), .ZN(\mexu/_0343_ ) );
XOR2_X1 \mexu/_1941_ ( .A(\mexu/_0199_ ), .B(\mexu/_1043_ ), .Z(\mexu/_0344_ ) );
INV_X1 \mexu/_1942_ ( .A(\mexu/_0344_ ), .ZN(\mexu/_0345_ ) );
OR2_X4 \mexu/_1943_ ( .A1(\mexu/_0343_ ), .A2(\mexu/_0345_ ), .ZN(\mexu/_0346_ ) );
AOI21_X1 \mexu/_1944_ ( .A(\mexu/_0794_ ), .B1(\mexu/_0343_ ), .B2(\mexu/_0345_ ), .ZN(\mexu/_0347_ ) );
NAND2_X1 \mexu/_1945_ ( .A1(\mexu/_0346_ ), .A2(\mexu/_0347_ ), .ZN(\mexu/_0348_ ) );
OR4_X4 \mexu/_1946_ ( .A1(\mexu/_0325_ ), .A2(\mexu/_0327_ ), .A3(\mexu/_0336_ ), .A4(\mexu/_0337_ ), .ZN(\mexu/_0349_ ) );
AOI21_X1 \mexu/_1947_ ( .A(\mexu/_0336_ ), .B1(\mexu/_0338_ ), .B2(\mexu/_0334_ ), .ZN(\mexu/_0350_ ) );
XOR2_X1 \mexu/_1948_ ( .A(\mexu/_0199_ ), .B(\mexu/_1001_ ), .Z(\mexu/_0351_ ) );
INV_X1 \mexu/_1949_ ( .A(\mexu/_0351_ ), .ZN(\mexu/_0352_ ) );
AND3_X2 \mexu/_1950_ ( .A1(\mexu/_0349_ ), .A2(\mexu/_0350_ ), .A3(\mexu/_0352_ ), .ZN(\mexu/_0353_ ) );
AOI21_X2 \mexu/_1951_ ( .A(\mexu/_0352_ ), .B1(\mexu/_0349_ ), .B2(\mexu/_0350_ ), .ZN(\mexu/_0354_ ) );
OR3_X2 \mexu/_1952_ ( .A1(\mexu/_0353_ ), .A2(\mexu/_0354_ ), .A3(\mexu/_0660_ ), .ZN(\mexu/_0355_ ) );
NAND2_X1 \mexu/_1953_ ( .A1(\mexu/_0348_ ), .A2(\mexu/_0355_ ), .ZN(\mexu/_0062_ ) );
NAND2_X1 \mexu/_1954_ ( .A1(\mexu/_0199_ ), .A2(\mexu/_1043_ ), .ZN(\mexu/_0356_ ) );
NAND2_X4 \mexu/_1955_ ( .A1(\mexu/_0346_ ), .A2(\mexu/_0356_ ), .ZN(\mexu/_0357_ ) );
XOR2_X1 \mexu/_1956_ ( .A(\mexu/_0200_ ), .B(\mexu/_1044_ ), .Z(\mexu/_0358_ ) );
AND2_X4 \mexu/_1957_ ( .A1(\mexu/_0357_ ), .A2(\mexu/_0358_ ), .ZN(\mexu/_0359_ ) );
OAI21_X1 \mexu/_1958_ ( .A(\mexu/_0661_ ), .B1(\mexu/_0357_ ), .B2(\mexu/_0358_ ), .ZN(\mexu/_0360_ ) );
AND2_X1 \mexu/_1959_ ( .A1(\mexu/_0199_ ), .A2(\mexu/_1001_ ), .ZN(\mexu/_0361_ ) );
NOR2_X1 \mexu/_1960_ ( .A1(\mexu/_0354_ ), .A2(\mexu/_0361_ ), .ZN(\mexu/_0362_ ) );
XNOR2_X1 \mexu/_1961_ ( .A(\mexu/_0200_ ), .B(\mexu/_1002_ ), .ZN(\mexu/_0363_ ) );
XNOR2_X2 \mexu/_1962_ ( .A(\mexu/_0362_ ), .B(\mexu/_0363_ ), .ZN(\mexu/_0364_ ) );
OAI22_X1 \mexu/_1963_ ( .A1(\mexu/_0359_ ), .A2(\mexu/_0360_ ), .B1(\mexu/_0776_ ), .B2(\mexu/_0364_ ), .ZN(\mexu/_0063_ ) );
NOR3_X1 \mexu/_1964_ ( .A1(\mexu/_0369_ ), .A2(\mexu/_0404_ ), .A3(\mexu/_0370_ ), .ZN(\mexu/_0209_ ) );
NOR3_X1 \mexu/_1965_ ( .A1(\mexu/_0369_ ), .A2(\mexu/_0406_ ), .A3(\mexu/_0370_ ), .ZN(\mexu/_0210_ ) );
NOR3_X1 \mexu/_1966_ ( .A1(\mexu/_0369_ ), .A2(\mexu/_0376_ ), .A3(\mexu/_0370_ ), .ZN(\mexu/_0211_ ) );
NOR3_X1 \mexu/_1967_ ( .A1(\mexu/_0369_ ), .A2(\mexu/_0378_ ), .A3(\mexu/_0402_ ), .ZN(\mexu/_0071_ ) );
AND3_X1 \mexu/_1968_ ( .A1(\mexu/_0213_ ), .A2(\mexu/_0434_ ), .A3(\mexu/_0437_ ), .ZN(\mexu/_0072_ ) );
AOI211_X4 \mexu/_1969_ ( .A(\mexu/_0175_ ), .B(\mexu/_0397_ ), .C1(\mexu/_0173_ ), .C2(\mexu/_0174_ ), .ZN(\mexu/_0172_ ) );
OAI211_X2 \mexu/_1970_ ( .A(\mexu/_0387_ ), .B(\mexu/_0380_ ), .C1(\mexu/_0973_ ), .C2(\mexu/_0365_ ), .ZN(\mexu/_0074_ ) );
DLL_X1 \mexu/_1971_ ( .D(\mexu/_1087_ ), .GN(upc_ctl ), .Q(\alu_ctl[0] ) );
DLL_X1 \mexu/_1972_ ( .D(\mexu/_1088_ ), .GN(upc_ctl ), .Q(\alu_ctl[1] ) );
DLL_X1 \mexu/_1973_ ( .D(\mexu/_1089_ ), .GN(upc_ctl ), .Q(\alu_ctl[2] ) );
DLL_X1 \mexu/_1974_ ( .D(\mexu/_1090_ ), .GN(upc_ctl ), .Q(\alu_ctl[3] ) );
DLL_X1 \mexu/_1975_ ( .D(mem_wen ), .GN(\mexu/_0036_ ), .Q(\wmask[0] ) );
DLL_X1 \mexu/_1976_ ( .D(\mexu/_0033_ ), .GN(\mexu/_0036_ ), .Q(\wmask[1] ) );
DLL_X1 \mexu/_1977_ ( .D(\mexu/_0035_ ), .GN(\mexu/_0036_ ), .Q(\wmask[3] ) );
DLH_X1 \mexu/_1978_ ( .D(\mexu/_1091_ ), .G(\mexu/_0038_ ), .Q(\csr_ctl[0] ) );
DLH_X1 \mexu/_1979_ ( .D(\mexu/_1092_ ), .G(\mexu/_0038_ ), .Q(\csr_ctl[1] ) );
DLH_X1 \mexu/_1980_ ( .D(\mexu/_1093_ ), .G(\mexu/_0038_ ), .Q(\csr_ctl[2] ) );
DLL_X1 \mexu/_1981_ ( .D(\mexu/_0000_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[0] ) );
DLL_X1 \mexu/_1982_ ( .D(\mexu/_0011_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[1] ) );
DLL_X1 \mexu/_1983_ ( .D(\mexu/_0022_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[2] ) );
DLL_X1 \mexu/_1984_ ( .D(\mexu/_0025_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[3] ) );
DLL_X1 \mexu/_1985_ ( .D(\mexu/_0026_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[4] ) );
DLL_X1 \mexu/_1986_ ( .D(\mexu/_0027_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[5] ) );
DLL_X1 \mexu/_1987_ ( .D(\mexu/_0028_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[6] ) );
DLL_X1 \mexu/_1988_ ( .D(\mexu/_0029_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[7] ) );
DLL_X1 \mexu/_1989_ ( .D(\mexu/_0030_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[8] ) );
DLL_X1 \mexu/_1990_ ( .D(\mexu/_0031_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[9] ) );
DLL_X1 \mexu/_1991_ ( .D(\mexu/_0001_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[10] ) );
DLL_X1 \mexu/_1992_ ( .D(\mexu/_0002_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[11] ) );
DLL_X1 \mexu/_1993_ ( .D(\mexu/_0003_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[12] ) );
DLL_X1 \mexu/_1994_ ( .D(\mexu/_0004_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[13] ) );
DLL_X1 \mexu/_1995_ ( .D(\mexu/_0005_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[14] ) );
DLL_X1 \mexu/_1996_ ( .D(\mexu/_0006_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[15] ) );
DLL_X1 \mexu/_1997_ ( .D(\mexu/_0007_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[16] ) );
DLL_X1 \mexu/_1998_ ( .D(\mexu/_0008_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[17] ) );
DLL_X1 \mexu/_1999_ ( .D(\mexu/_0009_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[18] ) );
DLL_X1 \mexu/_2000_ ( .D(\mexu/_0010_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[19] ) );
DLL_X1 \mexu/_2001_ ( .D(\mexu/_0012_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[20] ) );
DLL_X1 \mexu/_2002_ ( .D(\mexu/_0013_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[21] ) );
DLL_X1 \mexu/_2003_ ( .D(\mexu/_0014_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[22] ) );
DLL_X1 \mexu/_2004_ ( .D(\mexu/_0015_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[23] ) );
DLL_X1 \mexu/_2005_ ( .D(\mexu/_0016_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[24] ) );
DLL_X1 \mexu/_2006_ ( .D(\mexu/_0017_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[25] ) );
DLL_X1 \mexu/_2007_ ( .D(\mexu/_0018_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[26] ) );
DLL_X1 \mexu/_2008_ ( .D(\mexu/_0019_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[27] ) );
DLL_X1 \mexu/_2009_ ( .D(\mexu/_0020_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[28] ) );
DLL_X1 \mexu/_2010_ ( .D(\mexu/_0021_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[29] ) );
DLL_X1 \mexu/_2011_ ( .D(\mexu/_0023_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[30] ) );
DLL_X1 \mexu/_2012_ ( .D(\mexu/_0024_ ), .GN(\mexu/_0037_ ), .Q(\exu_upc[31] ) );
LOGIC0_X1 \mexu/_2013_ ( .Z(\mexu/_1086_ ) );
BUF_X1 \mexu/_2014_ ( .A(mem_wen ), .Z(\mexu/_0032_ ) );
BUF_X1 \mexu/_2015_ ( .A(\mexu/_0035_ ), .Z(\mexu/_0034_ ) );
BUF_X1 \mexu/_2016_ ( .A(mem_ren ), .Z(\result_ctl[0] ) );
BUF_X1 \mexu/_2017_ ( .A(\wmask[3] ), .Z(\wmask[2] ) );
BUF_X1 \mexu/_2018_ ( .A(\mexu/_1086_ ), .Z(\wmask[4] ) );
BUF_X1 \mexu/_2019_ ( .A(\mexu/_1086_ ), .Z(\wmask[5] ) );
BUF_X1 \mexu/_2020_ ( .A(\mexu/_1086_ ), .Z(\wmask[6] ) );
BUF_X1 \mexu/_2021_ ( .A(\mexu/_1086_ ), .Z(\wmask[7] ) );
BUF_X1 \mexu/_2022_ ( .A(\op[1] ), .Z(\mexu/_0972_ ) );
BUF_X1 \mexu/_2023_ ( .A(\op[0] ), .Z(\mexu/_0971_ ) );
BUF_X1 \mexu/_2024_ ( .A(\op[2] ), .Z(\mexu/_0973_ ) );
BUF_X1 \mexu/_2025_ ( .A(\op[3] ), .Z(\mexu/_0974_ ) );
BUF_X1 \mexu/_2026_ ( .A(\op[4] ), .Z(\mexu/_0975_ ) );
BUF_X1 \mexu/_2027_ ( .A(\op[5] ), .Z(\mexu/_0976_ ) );
BUF_X1 \mexu/_2028_ ( .A(\op[6] ), .Z(\mexu/_0977_ ) );
BUF_X1 \mexu/_2029_ ( .A(\mexu/_0212_ ), .Z(mem_ren ) );
BUF_X1 \mexu/_2030_ ( .A(\func[2] ), .Z(\mexu/_0175_ ) );
BUF_X1 \mexu/_2031_ ( .A(\func[0] ), .Z(\mexu/_0173_ ) );
BUF_X1 \mexu/_2032_ ( .A(\func[1] ), .Z(\mexu/_0174_ ) );
BUF_X1 \mexu/_2033_ ( .A(\mexu/_0075_ ), .Z(\mexu/_0038_ ) );
BUF_X1 \mexu/_2034_ ( .A(\mexu/_1085_ ), .Z(upc_ctl ) );
BUF_X1 \mexu/_2035_ ( .A(\mexu/_1017_ ), .Z(reg_wen ) );
BUF_X1 \mexu/_2036_ ( .A(\mexu/_0213_ ), .Z(mem_wen ) );
BUF_X1 \mexu/_2037_ ( .A(\mexu/_0073_ ), .Z(\mexu/_0036_ ) );
BUF_X1 \mexu/_2038_ ( .A(\imm[5] ), .Z(\mexu/_0203_ ) );
BUF_X1 \mexu/_2039_ ( .A(\imm[10] ), .Z(\mexu/_0177_ ) );
BUF_X1 \mexu/_2040_ ( .A(\mexu/_1010_ ), .Z(\mexu/_1087_ ) );
BUF_X1 \mexu/_2041_ ( .A(\mexu/_1011_ ), .Z(\mexu/_1088_ ) );
BUF_X1 \mexu/_2042_ ( .A(\mexu/_1012_ ), .Z(\mexu/_1089_ ) );
BUF_X1 \mexu/_2043_ ( .A(\mexu/_1013_ ), .Z(\mexu/_1090_ ) );
BUF_X1 \mexu/_2044_ ( .A(\imm[1] ), .Z(\mexu/_0187_ ) );
BUF_X1 \mexu/_2045_ ( .A(\imm[0] ), .Z(\mexu/_0176_ ) );
BUF_X1 \mexu/_2046_ ( .A(\mexu/_1014_ ), .Z(\mexu/_1091_ ) );
BUF_X1 \mexu/_2047_ ( .A(\mexu/_1015_ ), .Z(\mexu/_1092_ ) );
BUF_X1 \mexu/_2048_ ( .A(\mexu/_1016_ ), .Z(\mexu/_1093_ ) );
BUF_X1 \mexu/_2049_ ( .A(\csr_rdata[0] ), .Z(\mexu/_0140_ ) );
BUF_X1 \mexu/_2050_ ( .A(\mem_wdata[0] ), .Z(\mexu/_1052_ ) );
BUF_X1 \mexu/_2051_ ( .A(\mexu/_0108_ ), .Z(\alu_b[0] ) );
BUF_X1 \mexu/_2052_ ( .A(\csr_rdata[1] ), .Z(\mexu/_0151_ ) );
BUF_X1 \mexu/_2053_ ( .A(\mem_wdata[1] ), .Z(\mexu/_1063_ ) );
BUF_X1 \mexu/_2054_ ( .A(\mexu/_0119_ ), .Z(\alu_b[1] ) );
BUF_X1 \mexu/_2055_ ( .A(\csr_rdata[2] ), .Z(\mexu/_0162_ ) );
BUF_X1 \mexu/_2056_ ( .A(\mem_wdata[2] ), .Z(\mexu/_1074_ ) );
BUF_X1 \mexu/_2057_ ( .A(\imm[2] ), .Z(\mexu/_0198_ ) );
BUF_X1 \mexu/_2058_ ( .A(\mexu/_0130_ ), .Z(\alu_b[2] ) );
BUF_X1 \mexu/_2059_ ( .A(\csr_rdata[3] ), .Z(\mexu/_0165_ ) );
BUF_X1 \mexu/_2060_ ( .A(\mem_wdata[3] ), .Z(\mexu/_1077_ ) );
BUF_X1 \mexu/_2061_ ( .A(\imm[3] ), .Z(\mexu/_0201_ ) );
BUF_X1 \mexu/_2062_ ( .A(\mexu/_0133_ ), .Z(\alu_b[3] ) );
BUF_X1 \mexu/_2063_ ( .A(\csr_rdata[4] ), .Z(\mexu/_0166_ ) );
BUF_X1 \mexu/_2064_ ( .A(\mem_wdata[4] ), .Z(\mexu/_1078_ ) );
BUF_X1 \mexu/_2065_ ( .A(\imm[4] ), .Z(\mexu/_0202_ ) );
BUF_X1 \mexu/_2066_ ( .A(\mexu/_0134_ ), .Z(\alu_b[4] ) );
BUF_X1 \mexu/_2067_ ( .A(\csr_rdata[5] ), .Z(\mexu/_0167_ ) );
BUF_X1 \mexu/_2068_ ( .A(\mem_wdata[5] ), .Z(\mexu/_1079_ ) );
BUF_X1 \mexu/_2069_ ( .A(\mexu/_0135_ ), .Z(\alu_b[5] ) );
BUF_X1 \mexu/_2070_ ( .A(\csr_rdata[6] ), .Z(\mexu/_0168_ ) );
BUF_X1 \mexu/_2071_ ( .A(\mem_wdata[6] ), .Z(\mexu/_1080_ ) );
BUF_X1 \mexu/_2072_ ( .A(\imm[6] ), .Z(\mexu/_0204_ ) );
BUF_X1 \mexu/_2073_ ( .A(\mexu/_0136_ ), .Z(\alu_b[6] ) );
BUF_X1 \mexu/_2074_ ( .A(\csr_rdata[7] ), .Z(\mexu/_0169_ ) );
BUF_X1 \mexu/_2075_ ( .A(\mem_wdata[7] ), .Z(\mexu/_1081_ ) );
BUF_X1 \mexu/_2076_ ( .A(\imm[7] ), .Z(\mexu/_0205_ ) );
BUF_X1 \mexu/_2077_ ( .A(\mexu/_0137_ ), .Z(\alu_b[7] ) );
BUF_X1 \mexu/_2078_ ( .A(\csr_rdata[8] ), .Z(\mexu/_0170_ ) );
BUF_X1 \mexu/_2079_ ( .A(\mem_wdata[8] ), .Z(\mexu/_1082_ ) );
BUF_X1 \mexu/_2080_ ( .A(\imm[8] ), .Z(\mexu/_0206_ ) );
BUF_X1 \mexu/_2081_ ( .A(\mexu/_0138_ ), .Z(\alu_b[8] ) );
BUF_X1 \mexu/_2082_ ( .A(\csr_rdata[9] ), .Z(\mexu/_0171_ ) );
BUF_X1 \mexu/_2083_ ( .A(\mem_wdata[9] ), .Z(\mexu/_1083_ ) );
BUF_X1 \mexu/_2084_ ( .A(\imm[9] ), .Z(\mexu/_0207_ ) );
BUF_X1 \mexu/_2085_ ( .A(\mexu/_0139_ ), .Z(\alu_b[9] ) );
BUF_X1 \mexu/_2086_ ( .A(\csr_rdata[10] ), .Z(\mexu/_0141_ ) );
BUF_X1 \mexu/_2087_ ( .A(\mem_wdata[10] ), .Z(\mexu/_1053_ ) );
BUF_X1 \mexu/_2088_ ( .A(\mexu/_0109_ ), .Z(\alu_b[10] ) );
BUF_X1 \mexu/_2089_ ( .A(\csr_rdata[11] ), .Z(\mexu/_0142_ ) );
BUF_X1 \mexu/_2090_ ( .A(\mem_wdata[11] ), .Z(\mexu/_1054_ ) );
BUF_X1 \mexu/_2091_ ( .A(\imm[11] ), .Z(\mexu/_0178_ ) );
BUF_X1 \mexu/_2092_ ( .A(\mexu/_0110_ ), .Z(\alu_b[11] ) );
BUF_X1 \mexu/_2093_ ( .A(\csr_rdata[12] ), .Z(\mexu/_0143_ ) );
BUF_X1 \mexu/_2094_ ( .A(\mem_wdata[12] ), .Z(\mexu/_1055_ ) );
BUF_X1 \mexu/_2095_ ( .A(\imm[12] ), .Z(\mexu/_0179_ ) );
BUF_X1 \mexu/_2096_ ( .A(\mexu/_0111_ ), .Z(\alu_b[12] ) );
BUF_X1 \mexu/_2097_ ( .A(\csr_rdata[13] ), .Z(\mexu/_0144_ ) );
BUF_X1 \mexu/_2098_ ( .A(\mem_wdata[13] ), .Z(\mexu/_1056_ ) );
BUF_X1 \mexu/_2099_ ( .A(\imm[13] ), .Z(\mexu/_0180_ ) );
BUF_X1 \mexu/_2100_ ( .A(\mexu/_0112_ ), .Z(\alu_b[13] ) );
BUF_X1 \mexu/_2101_ ( .A(\csr_rdata[14] ), .Z(\mexu/_0145_ ) );
BUF_X1 \mexu/_2102_ ( .A(\mem_wdata[14] ), .Z(\mexu/_1057_ ) );
BUF_X1 \mexu/_2103_ ( .A(\imm[14] ), .Z(\mexu/_0181_ ) );
BUF_X1 \mexu/_2104_ ( .A(\mexu/_0113_ ), .Z(\alu_b[14] ) );
BUF_X1 \mexu/_2105_ ( .A(\csr_rdata[15] ), .Z(\mexu/_0146_ ) );
BUF_X1 \mexu/_2106_ ( .A(\mem_wdata[15] ), .Z(\mexu/_1058_ ) );
BUF_X1 \mexu/_2107_ ( .A(\imm[15] ), .Z(\mexu/_0182_ ) );
BUF_X1 \mexu/_2108_ ( .A(\mexu/_0114_ ), .Z(\alu_b[15] ) );
BUF_X1 \mexu/_2109_ ( .A(\csr_rdata[16] ), .Z(\mexu/_0147_ ) );
BUF_X1 \mexu/_2110_ ( .A(\mem_wdata[16] ), .Z(\mexu/_1059_ ) );
BUF_X1 \mexu/_2111_ ( .A(\imm[16] ), .Z(\mexu/_0183_ ) );
BUF_X1 \mexu/_2112_ ( .A(\mexu/_0115_ ), .Z(\alu_b[16] ) );
BUF_X1 \mexu/_2113_ ( .A(\csr_rdata[17] ), .Z(\mexu/_0148_ ) );
BUF_X1 \mexu/_2114_ ( .A(\mem_wdata[17] ), .Z(\mexu/_1060_ ) );
BUF_X1 \mexu/_2115_ ( .A(\imm[17] ), .Z(\mexu/_0184_ ) );
BUF_X1 \mexu/_2116_ ( .A(\mexu/_0116_ ), .Z(\alu_b[17] ) );
BUF_X1 \mexu/_2117_ ( .A(\csr_rdata[18] ), .Z(\mexu/_0149_ ) );
BUF_X1 \mexu/_2118_ ( .A(\mem_wdata[18] ), .Z(\mexu/_1061_ ) );
BUF_X1 \mexu/_2119_ ( .A(\imm[18] ), .Z(\mexu/_0185_ ) );
BUF_X1 \mexu/_2120_ ( .A(\mexu/_0117_ ), .Z(\alu_b[18] ) );
BUF_X1 \mexu/_2121_ ( .A(\csr_rdata[19] ), .Z(\mexu/_0150_ ) );
BUF_X1 \mexu/_2122_ ( .A(\mem_wdata[19] ), .Z(\mexu/_1062_ ) );
BUF_X1 \mexu/_2123_ ( .A(\imm[19] ), .Z(\mexu/_0186_ ) );
BUF_X1 \mexu/_2124_ ( .A(\mexu/_0118_ ), .Z(\alu_b[19] ) );
BUF_X1 \mexu/_2125_ ( .A(\csr_rdata[20] ), .Z(\mexu/_0152_ ) );
BUF_X1 \mexu/_2126_ ( .A(\mem_wdata[20] ), .Z(\mexu/_1064_ ) );
BUF_X1 \mexu/_2127_ ( .A(\imm[20] ), .Z(\mexu/_0188_ ) );
BUF_X1 \mexu/_2128_ ( .A(\mexu/_0120_ ), .Z(\alu_b[20] ) );
BUF_X1 \mexu/_2129_ ( .A(\csr_rdata[21] ), .Z(\mexu/_0153_ ) );
BUF_X1 \mexu/_2130_ ( .A(\mem_wdata[21] ), .Z(\mexu/_1065_ ) );
BUF_X1 \mexu/_2131_ ( .A(\imm[21] ), .Z(\mexu/_0189_ ) );
BUF_X1 \mexu/_2132_ ( .A(\mexu/_0121_ ), .Z(\alu_b[21] ) );
BUF_X1 \mexu/_2133_ ( .A(\csr_rdata[22] ), .Z(\mexu/_0154_ ) );
BUF_X1 \mexu/_2134_ ( .A(\mem_wdata[22] ), .Z(\mexu/_1066_ ) );
BUF_X1 \mexu/_2135_ ( .A(\imm[22] ), .Z(\mexu/_0190_ ) );
BUF_X1 \mexu/_2136_ ( .A(\mexu/_0122_ ), .Z(\alu_b[22] ) );
BUF_X1 \mexu/_2137_ ( .A(\csr_rdata[23] ), .Z(\mexu/_0155_ ) );
BUF_X1 \mexu/_2138_ ( .A(\mem_wdata[23] ), .Z(\mexu/_1067_ ) );
BUF_X1 \mexu/_2139_ ( .A(\imm[23] ), .Z(\mexu/_0191_ ) );
BUF_X1 \mexu/_2140_ ( .A(\mexu/_0123_ ), .Z(\alu_b[23] ) );
BUF_X1 \mexu/_2141_ ( .A(\csr_rdata[24] ), .Z(\mexu/_0156_ ) );
BUF_X1 \mexu/_2142_ ( .A(\mem_wdata[24] ), .Z(\mexu/_1068_ ) );
BUF_X1 \mexu/_2143_ ( .A(\imm[24] ), .Z(\mexu/_0192_ ) );
BUF_X1 \mexu/_2144_ ( .A(\mexu/_0124_ ), .Z(\alu_b[24] ) );
BUF_X1 \mexu/_2145_ ( .A(\csr_rdata[25] ), .Z(\mexu/_0157_ ) );
BUF_X1 \mexu/_2146_ ( .A(\mem_wdata[25] ), .Z(\mexu/_1069_ ) );
BUF_X1 \mexu/_2147_ ( .A(\imm[25] ), .Z(\mexu/_0193_ ) );
BUF_X1 \mexu/_2148_ ( .A(\mexu/_0125_ ), .Z(\alu_b[25] ) );
BUF_X1 \mexu/_2149_ ( .A(\csr_rdata[26] ), .Z(\mexu/_0158_ ) );
BUF_X1 \mexu/_2150_ ( .A(\mem_wdata[26] ), .Z(\mexu/_1070_ ) );
BUF_X1 \mexu/_2151_ ( .A(\imm[26] ), .Z(\mexu/_0194_ ) );
BUF_X1 \mexu/_2152_ ( .A(\mexu/_0126_ ), .Z(\alu_b[26] ) );
BUF_X1 \mexu/_2153_ ( .A(\csr_rdata[27] ), .Z(\mexu/_0159_ ) );
BUF_X1 \mexu/_2154_ ( .A(\mem_wdata[27] ), .Z(\mexu/_1071_ ) );
BUF_X1 \mexu/_2155_ ( .A(\imm[27] ), .Z(\mexu/_0195_ ) );
BUF_X1 \mexu/_2156_ ( .A(\mexu/_0127_ ), .Z(\alu_b[27] ) );
BUF_X1 \mexu/_2157_ ( .A(\csr_rdata[28] ), .Z(\mexu/_0160_ ) );
BUF_X1 \mexu/_2158_ ( .A(\mem_wdata[28] ), .Z(\mexu/_1072_ ) );
BUF_X1 \mexu/_2159_ ( .A(\imm[28] ), .Z(\mexu/_0196_ ) );
BUF_X1 \mexu/_2160_ ( .A(\mexu/_0128_ ), .Z(\alu_b[28] ) );
BUF_X1 \mexu/_2161_ ( .A(\csr_rdata[29] ), .Z(\mexu/_0161_ ) );
BUF_X1 \mexu/_2162_ ( .A(\mem_wdata[29] ), .Z(\mexu/_1073_ ) );
BUF_X1 \mexu/_2163_ ( .A(\imm[29] ), .Z(\mexu/_0197_ ) );
BUF_X1 \mexu/_2164_ ( .A(\mexu/_0129_ ), .Z(\alu_b[29] ) );
BUF_X1 \mexu/_2165_ ( .A(\csr_rdata[30] ), .Z(\mexu/_0163_ ) );
BUF_X1 \mexu/_2166_ ( .A(\mem_wdata[30] ), .Z(\mexu/_1075_ ) );
BUF_X1 \mexu/_2167_ ( .A(\imm[30] ), .Z(\mexu/_0199_ ) );
BUF_X1 \mexu/_2168_ ( .A(\mexu/_0131_ ), .Z(\alu_b[30] ) );
BUF_X1 \mexu/_2169_ ( .A(\csr_rdata[31] ), .Z(\mexu/_0164_ ) );
BUF_X1 \mexu/_2170_ ( .A(\mem_wdata[31] ), .Z(\mexu/_1076_ ) );
BUF_X1 \mexu/_2171_ ( .A(\imm[31] ), .Z(\mexu/_0200_ ) );
BUF_X1 \mexu/_2172_ ( .A(\mexu/_0132_ ), .Z(\alu_b[31] ) );
BUF_X1 \mexu/_2173_ ( .A(\pc[0] ), .Z(\mexu/_0978_ ) );
BUF_X1 \mexu/_2174_ ( .A(\src1[0] ), .Z(\mexu/_1020_ ) );
BUF_X1 \mexu/_2175_ ( .A(\mexu/_0076_ ), .Z(\alu_a[0] ) );
BUF_X1 \mexu/_2176_ ( .A(\pc[1] ), .Z(\mexu/_0989_ ) );
BUF_X1 \mexu/_2177_ ( .A(\src1[1] ), .Z(\mexu/_1031_ ) );
BUF_X1 \mexu/_2178_ ( .A(\mexu/_0087_ ), .Z(\alu_a[1] ) );
BUF_X1 \mexu/_2179_ ( .A(\pc[2] ), .Z(\mexu/_1000_ ) );
BUF_X1 \mexu/_2180_ ( .A(\src1[2] ), .Z(\mexu/_1042_ ) );
BUF_X1 \mexu/_2181_ ( .A(\mexu/_0098_ ), .Z(\alu_a[2] ) );
BUF_X1 \mexu/_2182_ ( .A(\pc[3] ), .Z(\mexu/_1003_ ) );
BUF_X1 \mexu/_2183_ ( .A(\src1[3] ), .Z(\mexu/_1045_ ) );
BUF_X1 \mexu/_2184_ ( .A(\mexu/_0101_ ), .Z(\alu_a[3] ) );
BUF_X1 \mexu/_2185_ ( .A(\pc[4] ), .Z(\mexu/_1004_ ) );
BUF_X1 \mexu/_2186_ ( .A(\src1[4] ), .Z(\mexu/_1046_ ) );
BUF_X1 \mexu/_2187_ ( .A(\mexu/_0102_ ), .Z(\alu_a[4] ) );
BUF_X1 \mexu/_2188_ ( .A(\pc[5] ), .Z(\mexu/_1005_ ) );
BUF_X1 \mexu/_2189_ ( .A(\src1[5] ), .Z(\mexu/_1047_ ) );
BUF_X1 \mexu/_2190_ ( .A(\mexu/_0103_ ), .Z(\alu_a[5] ) );
BUF_X1 \mexu/_2191_ ( .A(\pc[6] ), .Z(\mexu/_1006_ ) );
BUF_X1 \mexu/_2192_ ( .A(\src1[6] ), .Z(\mexu/_1048_ ) );
BUF_X1 \mexu/_2193_ ( .A(\mexu/_0104_ ), .Z(\alu_a[6] ) );
BUF_X1 \mexu/_2194_ ( .A(\pc[7] ), .Z(\mexu/_1007_ ) );
BUF_X1 \mexu/_2195_ ( .A(\src1[7] ), .Z(\mexu/_1049_ ) );
BUF_X1 \mexu/_2196_ ( .A(\mexu/_0105_ ), .Z(\alu_a[7] ) );
BUF_X1 \mexu/_2197_ ( .A(\pc[8] ), .Z(\mexu/_1008_ ) );
BUF_X1 \mexu/_2198_ ( .A(\src1[8] ), .Z(\mexu/_1050_ ) );
BUF_X1 \mexu/_2199_ ( .A(\mexu/_0106_ ), .Z(\alu_a[8] ) );
BUF_X1 \mexu/_2200_ ( .A(\pc[9] ), .Z(\mexu/_1009_ ) );
BUF_X1 \mexu/_2201_ ( .A(\src1[9] ), .Z(\mexu/_1051_ ) );
BUF_X1 \mexu/_2202_ ( .A(\mexu/_0107_ ), .Z(\alu_a[9] ) );
BUF_X1 \mexu/_2203_ ( .A(\pc[10] ), .Z(\mexu/_0979_ ) );
BUF_X1 \mexu/_2204_ ( .A(\src1[10] ), .Z(\mexu/_1021_ ) );
BUF_X1 \mexu/_2205_ ( .A(\mexu/_0077_ ), .Z(\alu_a[10] ) );
BUF_X1 \mexu/_2206_ ( .A(\pc[11] ), .Z(\mexu/_0980_ ) );
BUF_X1 \mexu/_2207_ ( .A(\src1[11] ), .Z(\mexu/_1022_ ) );
BUF_X1 \mexu/_2208_ ( .A(\mexu/_0078_ ), .Z(\alu_a[11] ) );
BUF_X1 \mexu/_2209_ ( .A(\pc[12] ), .Z(\mexu/_0981_ ) );
BUF_X1 \mexu/_2210_ ( .A(\src1[12] ), .Z(\mexu/_1023_ ) );
BUF_X1 \mexu/_2211_ ( .A(\mexu/_0079_ ), .Z(\alu_a[12] ) );
BUF_X1 \mexu/_2212_ ( .A(\pc[13] ), .Z(\mexu/_0982_ ) );
BUF_X1 \mexu/_2213_ ( .A(\src1[13] ), .Z(\mexu/_1024_ ) );
BUF_X1 \mexu/_2214_ ( .A(\mexu/_0080_ ), .Z(\alu_a[13] ) );
BUF_X1 \mexu/_2215_ ( .A(\pc[14] ), .Z(\mexu/_0983_ ) );
BUF_X1 \mexu/_2216_ ( .A(\src1[14] ), .Z(\mexu/_1025_ ) );
BUF_X1 \mexu/_2217_ ( .A(\mexu/_0081_ ), .Z(\alu_a[14] ) );
BUF_X1 \mexu/_2218_ ( .A(\pc[15] ), .Z(\mexu/_0984_ ) );
BUF_X1 \mexu/_2219_ ( .A(\src1[15] ), .Z(\mexu/_1026_ ) );
BUF_X1 \mexu/_2220_ ( .A(\mexu/_0082_ ), .Z(\alu_a[15] ) );
BUF_X1 \mexu/_2221_ ( .A(\pc[16] ), .Z(\mexu/_0985_ ) );
BUF_X1 \mexu/_2222_ ( .A(\src1[16] ), .Z(\mexu/_1027_ ) );
BUF_X1 \mexu/_2223_ ( .A(\mexu/_0083_ ), .Z(\alu_a[16] ) );
BUF_X1 \mexu/_2224_ ( .A(\pc[17] ), .Z(\mexu/_0986_ ) );
BUF_X1 \mexu/_2225_ ( .A(\src1[17] ), .Z(\mexu/_1028_ ) );
BUF_X1 \mexu/_2226_ ( .A(\mexu/_0084_ ), .Z(\alu_a[17] ) );
BUF_X1 \mexu/_2227_ ( .A(\pc[18] ), .Z(\mexu/_0987_ ) );
BUF_X1 \mexu/_2228_ ( .A(\src1[18] ), .Z(\mexu/_1029_ ) );
BUF_X1 \mexu/_2229_ ( .A(\mexu/_0085_ ), .Z(\alu_a[18] ) );
BUF_X1 \mexu/_2230_ ( .A(\pc[19] ), .Z(\mexu/_0988_ ) );
BUF_X1 \mexu/_2231_ ( .A(\src1[19] ), .Z(\mexu/_1030_ ) );
BUF_X1 \mexu/_2232_ ( .A(\mexu/_0086_ ), .Z(\alu_a[19] ) );
BUF_X1 \mexu/_2233_ ( .A(\pc[20] ), .Z(\mexu/_0990_ ) );
BUF_X1 \mexu/_2234_ ( .A(\src1[20] ), .Z(\mexu/_1032_ ) );
BUF_X1 \mexu/_2235_ ( .A(\mexu/_0088_ ), .Z(\alu_a[20] ) );
BUF_X1 \mexu/_2236_ ( .A(\pc[21] ), .Z(\mexu/_0991_ ) );
BUF_X1 \mexu/_2237_ ( .A(\src1[21] ), .Z(\mexu/_1033_ ) );
BUF_X1 \mexu/_2238_ ( .A(\mexu/_0089_ ), .Z(\alu_a[21] ) );
BUF_X1 \mexu/_2239_ ( .A(\pc[22] ), .Z(\mexu/_0992_ ) );
BUF_X1 \mexu/_2240_ ( .A(\src1[22] ), .Z(\mexu/_1034_ ) );
BUF_X1 \mexu/_2241_ ( .A(\mexu/_0090_ ), .Z(\alu_a[22] ) );
BUF_X1 \mexu/_2242_ ( .A(\pc[23] ), .Z(\mexu/_0993_ ) );
BUF_X1 \mexu/_2243_ ( .A(\src1[23] ), .Z(\mexu/_1035_ ) );
BUF_X1 \mexu/_2244_ ( .A(\mexu/_0091_ ), .Z(\alu_a[23] ) );
BUF_X1 \mexu/_2245_ ( .A(\pc[24] ), .Z(\mexu/_0994_ ) );
BUF_X1 \mexu/_2246_ ( .A(\src1[24] ), .Z(\mexu/_1036_ ) );
BUF_X1 \mexu/_2247_ ( .A(\mexu/_0092_ ), .Z(\alu_a[24] ) );
BUF_X1 \mexu/_2248_ ( .A(\pc[25] ), .Z(\mexu/_0995_ ) );
BUF_X1 \mexu/_2249_ ( .A(\src1[25] ), .Z(\mexu/_1037_ ) );
BUF_X1 \mexu/_2250_ ( .A(\mexu/_0093_ ), .Z(\alu_a[25] ) );
BUF_X1 \mexu/_2251_ ( .A(\pc[26] ), .Z(\mexu/_0996_ ) );
BUF_X1 \mexu/_2252_ ( .A(\src1[26] ), .Z(\mexu/_1038_ ) );
BUF_X1 \mexu/_2253_ ( .A(\mexu/_0094_ ), .Z(\alu_a[26] ) );
BUF_X1 \mexu/_2254_ ( .A(\pc[27] ), .Z(\mexu/_0997_ ) );
BUF_X1 \mexu/_2255_ ( .A(\src1[27] ), .Z(\mexu/_1039_ ) );
BUF_X1 \mexu/_2256_ ( .A(\mexu/_0095_ ), .Z(\alu_a[27] ) );
BUF_X1 \mexu/_2257_ ( .A(\pc[28] ), .Z(\mexu/_0998_ ) );
BUF_X1 \mexu/_2258_ ( .A(\src1[28] ), .Z(\mexu/_1040_ ) );
BUF_X1 \mexu/_2259_ ( .A(\mexu/_0096_ ), .Z(\alu_a[28] ) );
BUF_X1 \mexu/_2260_ ( .A(\pc[29] ), .Z(\mexu/_0999_ ) );
BUF_X1 \mexu/_2261_ ( .A(\src1[29] ), .Z(\mexu/_1041_ ) );
BUF_X1 \mexu/_2262_ ( .A(\mexu/_0097_ ), .Z(\alu_a[29] ) );
BUF_X1 \mexu/_2263_ ( .A(\pc[30] ), .Z(\mexu/_1001_ ) );
BUF_X1 \mexu/_2264_ ( .A(\src1[30] ), .Z(\mexu/_1043_ ) );
BUF_X1 \mexu/_2265_ ( .A(\mexu/_0099_ ), .Z(\alu_a[30] ) );
BUF_X1 \mexu/_2266_ ( .A(\pc[31] ), .Z(\mexu/_1002_ ) );
BUF_X1 \mexu/_2267_ ( .A(\src1[31] ), .Z(\mexu/_1044_ ) );
BUF_X1 \mexu/_2268_ ( .A(\mexu/_0100_ ), .Z(\alu_a[31] ) );
BUF_X1 \mexu/_2269_ ( .A(\mexu/_1019_ ), .Z(alu_sign ) );
BUF_X1 \mexu/_2270_ ( .A(\mexu/_1084_ ), .Z(alu_sub ) );
BUF_X1 \mexu/_2271_ ( .A(\mexu/_1018_ ), .Z(\result_ctl[1] ) );
BUF_X1 \mexu/_2272_ ( .A(\mexu/_0208_ ), .Z(exu_jump ) );
BUF_X1 \mexu/_2273_ ( .A(\mexu/_0039_ ), .Z(\mexu/_0000_ ) );
BUF_X1 \mexu/_2274_ ( .A(\mexu/_0050_ ), .Z(\mexu/_0011_ ) );
BUF_X1 \mexu/_2275_ ( .A(\mexu/_0061_ ), .Z(\mexu/_0022_ ) );
BUF_X1 \mexu/_2276_ ( .A(\mexu/_0064_ ), .Z(\mexu/_0025_ ) );
BUF_X1 \mexu/_2277_ ( .A(\mexu/_0065_ ), .Z(\mexu/_0026_ ) );
BUF_X1 \mexu/_2278_ ( .A(\mexu/_0066_ ), .Z(\mexu/_0027_ ) );
BUF_X1 \mexu/_2279_ ( .A(\mexu/_0067_ ), .Z(\mexu/_0028_ ) );
BUF_X1 \mexu/_2280_ ( .A(\mexu/_0068_ ), .Z(\mexu/_0029_ ) );
BUF_X1 \mexu/_2281_ ( .A(\mexu/_0069_ ), .Z(\mexu/_0030_ ) );
BUF_X1 \mexu/_2282_ ( .A(\mexu/_0070_ ), .Z(\mexu/_0031_ ) );
BUF_X1 \mexu/_2283_ ( .A(\mexu/_0040_ ), .Z(\mexu/_0001_ ) );
BUF_X1 \mexu/_2284_ ( .A(\mexu/_0041_ ), .Z(\mexu/_0002_ ) );
BUF_X1 \mexu/_2285_ ( .A(\mexu/_0042_ ), .Z(\mexu/_0003_ ) );
BUF_X1 \mexu/_2286_ ( .A(\mexu/_0043_ ), .Z(\mexu/_0004_ ) );
BUF_X1 \mexu/_2287_ ( .A(\mexu/_0044_ ), .Z(\mexu/_0005_ ) );
BUF_X1 \mexu/_2288_ ( .A(\mexu/_0045_ ), .Z(\mexu/_0006_ ) );
BUF_X1 \mexu/_2289_ ( .A(\mexu/_0046_ ), .Z(\mexu/_0007_ ) );
BUF_X1 \mexu/_2290_ ( .A(\mexu/_0047_ ), .Z(\mexu/_0008_ ) );
BUF_X1 \mexu/_2291_ ( .A(\mexu/_0048_ ), .Z(\mexu/_0009_ ) );
BUF_X1 \mexu/_2292_ ( .A(\mexu/_0049_ ), .Z(\mexu/_0010_ ) );
BUF_X1 \mexu/_2293_ ( .A(\mexu/_0051_ ), .Z(\mexu/_0012_ ) );
BUF_X1 \mexu/_2294_ ( .A(\mexu/_0052_ ), .Z(\mexu/_0013_ ) );
BUF_X1 \mexu/_2295_ ( .A(\mexu/_0053_ ), .Z(\mexu/_0014_ ) );
BUF_X1 \mexu/_2296_ ( .A(\mexu/_0054_ ), .Z(\mexu/_0015_ ) );
BUF_X1 \mexu/_2297_ ( .A(\mexu/_0055_ ), .Z(\mexu/_0016_ ) );
BUF_X1 \mexu/_2298_ ( .A(\mexu/_0056_ ), .Z(\mexu/_0017_ ) );
BUF_X1 \mexu/_2299_ ( .A(\mexu/_0057_ ), .Z(\mexu/_0018_ ) );
BUF_X1 \mexu/_2300_ ( .A(\mexu/_0058_ ), .Z(\mexu/_0019_ ) );
BUF_X1 \mexu/_2301_ ( .A(\mexu/_0059_ ), .Z(\mexu/_0020_ ) );
BUF_X1 \mexu/_2302_ ( .A(\mexu/_0060_ ), .Z(\mexu/_0021_ ) );
BUF_X1 \mexu/_2303_ ( .A(\mexu/_0062_ ), .Z(\mexu/_0023_ ) );
BUF_X1 \mexu/_2304_ ( .A(\mexu/_0063_ ), .Z(\mexu/_0024_ ) );
BUF_X1 \mexu/_2305_ ( .A(\mexu/_0209_ ), .Z(\load_ctl[0] ) );
BUF_X1 \mexu/_2306_ ( .A(\mexu/_0210_ ), .Z(\load_ctl[1] ) );
BUF_X1 \mexu/_2307_ ( .A(\mexu/_0211_ ), .Z(\load_ctl[2] ) );
BUF_X1 \mexu/_2308_ ( .A(\mexu/_0071_ ), .Z(\mexu/_0033_ ) );
BUF_X1 \mexu/_2309_ ( .A(\mexu/_0072_ ), .Z(\mexu/_0035_ ) );
BUF_X1 \mexu/_2310_ ( .A(\mexu/_0172_ ), .Z(csr_wen ) );
BUF_X1 \mexu/_2311_ ( .A(\mexu/_0074_ ), .Z(\mexu/_0037_ ) );
AND2_X4 \midu/_131_ ( .A1(\midu/_043_ ), .A2(\midu/_032_ ), .ZN(\midu/_098_ ) );
NOR2_X4 \midu/_132_ ( .A1(\midu/_057_ ), .A2(\midu/_054_ ), .ZN(\midu/_099_ ) );
AND2_X4 \midu/_133_ ( .A1(\midu/_098_ ), .A2(\midu/_099_ ), .ZN(\midu/_100_ ) );
INV_X32 \midu/_134_ ( .A(\midu/_059_ ), .ZN(\midu/_101_ ) );
NOR2_X4 \midu/_135_ ( .A1(\midu/_101_ ), .A2(\midu/_058_ ), .ZN(\midu/_102_ ) );
AND2_X2 \midu/_136_ ( .A1(\midu/_100_ ), .A2(\midu/_102_ ), .ZN(\midu/_103_ ) );
INV_X1 \midu/_137_ ( .A(\midu/_060_ ), .ZN(\midu/_104_ ) );
NAND3_X1 \midu/_138_ ( .A1(\midu/_103_ ), .A2(\midu/_104_ ), .A3(\midu/_061_ ), .ZN(\midu/_105_ ) );
AND3_X1 \midu/_139_ ( .A1(\midu/_104_ ), .A2(\midu/_059_ ), .A3(\midu/_058_ ), .ZN(\midu/_106_ ) );
AND2_X1 \midu/_140_ ( .A1(\midu/_100_ ), .A2(\midu/_106_ ), .ZN(\midu/_107_ ) );
INV_X1 \midu/_141_ ( .A(\midu/_107_ ), .ZN(\midu/_108_ ) );
INV_X1 \midu/_142_ ( .A(\midu/_049_ ), .ZN(\midu/_109_ ) );
INV_X1 \midu/_143_ ( .A(\midu/_058_ ), .ZN(\midu/_110_ ) );
NAND4_X2 \midu/_144_ ( .A1(\midu/_100_ ), .A2(\midu/_101_ ), .A3(\midu/_110_ ), .A4(\midu/_104_ ), .ZN(\midu/_111_ ) );
NAND4_X2 \midu/_145_ ( .A1(\midu/_100_ ), .A2(\midu/_101_ ), .A3(\midu/_058_ ), .A4(\midu/_104_ ), .ZN(\midu/_112_ ) );
NAND2_X2 \midu/_146_ ( .A1(\midu/_111_ ), .A2(\midu/_112_ ), .ZN(\midu/_113_ ) );
NAND3_X1 \midu/_147_ ( .A1(\midu/_043_ ), .A2(\midu/_032_ ), .A3(\midu/_054_ ), .ZN(\midu/_114_ ) );
NOR2_X1 \midu/_148_ ( .A1(\midu/_114_ ), .A2(\midu/_057_ ), .ZN(\midu/_115_ ) );
NAND3_X1 \midu/_149_ ( .A1(\midu/_115_ ), .A2(\midu/_060_ ), .A3(\midu/_102_ ), .ZN(\midu/_116_ ) );
AND2_X2 \midu/_150_ ( .A1(\midu/_059_ ), .A2(\midu/_058_ ), .ZN(\midu/_117_ ) );
NAND4_X1 \midu/_151_ ( .A1(\midu/_098_ ), .A2(\midu/_117_ ), .A3(\midu/_060_ ), .A4(\midu/_099_ ), .ZN(\midu/_118_ ) );
NAND2_X4 \midu/_152_ ( .A1(\midu/_116_ ), .A2(\midu/_118_ ), .ZN(\midu/_119_ ) );
NOR2_X4 \midu/_153_ ( .A1(\midu/_113_ ), .A2(\midu/_119_ ), .ZN(\midu/_120_ ) );
INV_X1 \midu/_154_ ( .A(\midu/_044_ ), .ZN(\midu/_121_ ) );
OAI221_X1 \midu/_155_ ( .A(\midu/_105_ ), .B1(\midu/_108_ ), .B2(\midu/_109_ ), .C1(\midu/_120_ ), .C2(\midu/_121_ ), .ZN(\midu/_000_ ) );
NAND4_X1 \midu/_156_ ( .A1(\midu/_102_ ), .A2(\midu/_062_ ), .A3(\midu/_098_ ), .A4(\midu/_099_ ), .ZN(\midu/_122_ ) );
INV_X1 \midu/_157_ ( .A(\midu/_050_ ), .ZN(\midu/_123_ ) );
AND2_X4 \midu/_158_ ( .A1(\midu/_102_ ), .A2(\midu/_060_ ), .ZN(\midu/_124_ ) );
AND4_X4 \midu/_159_ ( .A1(\midu/_043_ ), .A2(\midu/_032_ ), .A3(\midu/_057_ ), .A4(\midu/_054_ ), .ZN(\midu/_125_ ) );
AND2_X4 \midu/_160_ ( .A1(\midu/_124_ ), .A2(\midu/_125_ ), .ZN(\midu/_126_ ) );
BUF_X8 \midu/_161_ ( .A(\midu/_126_ ), .Z(\midu/_127_ ) );
INV_X1 \midu/_162_ ( .A(\midu/_127_ ), .ZN(\midu/_128_ ) );
AND2_X4 \midu/_163_ ( .A1(\midu/_120_ ), .A2(\midu/_128_ ), .ZN(\midu/_129_ ) );
INV_X1 \midu/_164_ ( .A(\midu/_045_ ), .ZN(\midu/_130_ ) );
OAI221_X1 \midu/_165_ ( .A(\midu/_122_ ), .B1(\midu/_123_ ), .B2(\midu/_108_ ), .C1(\midu/_129_ ), .C2(\midu/_130_ ), .ZN(\midu/_011_ ) );
NAND4_X1 \midu/_166_ ( .A1(\midu/_102_ ), .A2(\midu/_063_ ), .A3(\midu/_098_ ), .A4(\midu/_099_ ), .ZN(\midu/_064_ ) );
INV_X1 \midu/_167_ ( .A(\midu/_051_ ), .ZN(\midu/_065_ ) );
INV_X1 \midu/_168_ ( .A(\midu/_046_ ), .ZN(\midu/_066_ ) );
OAI221_X1 \midu/_169_ ( .A(\midu/_064_ ), .B1(\midu/_065_ ), .B2(\midu/_108_ ), .C1(\midu/_129_ ), .C2(\midu/_066_ ), .ZN(\midu/_022_ ) );
NAND4_X1 \midu/_170_ ( .A1(\midu/_102_ ), .A2(\midu/_033_ ), .A3(\midu/_098_ ), .A4(\midu/_099_ ), .ZN(\midu/_067_ ) );
INV_X1 \midu/_171_ ( .A(\midu/_052_ ), .ZN(\midu/_068_ ) );
INV_X1 \midu/_172_ ( .A(\midu/_047_ ), .ZN(\midu/_069_ ) );
OAI221_X1 \midu/_173_ ( .A(\midu/_067_ ), .B1(\midu/_068_ ), .B2(\midu/_108_ ), .C1(\midu/_129_ ), .C2(\midu/_069_ ), .ZN(\midu/_025_ ) );
NAND4_X1 \midu/_174_ ( .A1(\midu/_102_ ), .A2(\midu/_034_ ), .A3(\midu/_098_ ), .A4(\midu/_099_ ), .ZN(\midu/_070_ ) );
INV_X1 \midu/_175_ ( .A(\midu/_053_ ), .ZN(\midu/_071_ ) );
INV_X1 \midu/_176_ ( .A(\midu/_048_ ), .ZN(\midu/_072_ ) );
OAI221_X1 \midu/_177_ ( .A(\midu/_070_ ), .B1(\midu/_071_ ), .B2(\midu/_108_ ), .C1(\midu/_129_ ), .C2(\midu/_072_ ), .ZN(\midu/_026_ ) );
NOR2_X2 \midu/_178_ ( .A1(\midu/_127_ ), .A2(\midu/_103_ ), .ZN(\midu/_073_ ) );
AND2_X4 \midu/_179_ ( .A1(\midu/_120_ ), .A2(\midu/_073_ ), .ZN(\midu/_074_ ) );
BUF_X8 \midu/_180_ ( .A(\midu/_074_ ), .Z(\midu/_075_ ) );
INV_X1 \midu/_181_ ( .A(\midu/_055_ ), .ZN(\midu/_076_ ) );
OAI22_X1 \midu/_182_ ( .A1(\midu/_075_ ), .A2(\midu/_109_ ), .B1(\midu/_076_ ), .B2(\midu/_108_ ), .ZN(\midu/_027_ ) );
INV_X1 \midu/_183_ ( .A(\midu/_056_ ), .ZN(\midu/_077_ ) );
OAI22_X1 \midu/_184_ ( .A1(\midu/_075_ ), .A2(\midu/_123_ ), .B1(\midu/_077_ ), .B2(\midu/_108_ ), .ZN(\midu/_028_ ) );
AOI21_X1 \midu/_185_ ( .A(\midu/_065_ ), .B1(\midu/_120_ ), .B2(\midu/_073_ ), .ZN(\midu/_029_ ) );
AOI21_X1 \midu/_186_ ( .A(\midu/_068_ ), .B1(\midu/_120_ ), .B2(\midu/_073_ ), .ZN(\midu/_030_ ) );
AOI21_X1 \midu/_187_ ( .A(\midu/_071_ ), .B1(\midu/_120_ ), .B2(\midu/_073_ ), .ZN(\midu/_031_ ) );
AOI21_X1 \midu/_188_ ( .A(\midu/_076_ ), .B1(\midu/_120_ ), .B2(\midu/_073_ ), .ZN(\midu/_001_ ) );
AND3_X1 \midu/_189_ ( .A1(\midu/_124_ ), .A2(\midu/_061_ ), .A3(\midu/_100_ ), .ZN(\midu/_078_ ) );
AND2_X1 \midu/_190_ ( .A1(\midu/_103_ ), .A2(\midu/_104_ ), .ZN(\midu/_079_ ) );
AOI21_X1 \midu/_191_ ( .A(\midu/_078_ ), .B1(\midu/_079_ ), .B2(\midu/_056_ ), .ZN(\midu/_080_ ) );
OAI221_X1 \midu/_192_ ( .A(\midu/_080_ ), .B1(\midu/_121_ ), .B2(\midu/_128_ ), .C1(\midu/_077_ ), .C2(\midu/_120_ ), .ZN(\midu/_002_ ) );
NOR2_X2 \midu/_193_ ( .A1(\midu/_120_ ), .A2(\midu/_077_ ), .ZN(\midu/_081_ ) );
AND4_X1 \midu/_194_ ( .A1(\midu/_056_ ), .A2(\midu/_102_ ), .A3(\midu/_098_ ), .A4(\midu/_099_ ), .ZN(\midu/_082_ ) );
NOR2_X4 \midu/_195_ ( .A1(\midu/_081_ ), .A2(\midu/_082_ ), .ZN(\midu/_083_ ) );
NOR2_X1 \midu/_196_ ( .A1(\midu/_110_ ), .A2(\midu/_060_ ), .ZN(\midu/_084_ ) );
AND2_X2 \midu/_197_ ( .A1(\midu/_115_ ), .A2(\midu/_084_ ), .ZN(\midu/_085_ ) );
OAI21_X1 \midu/_198_ ( .A(\midu/_035_ ), .B1(\midu/_127_ ), .B2(\midu/_085_ ), .ZN(\midu/_086_ ) );
NAND2_X1 \midu/_199_ ( .A1(\midu/_083_ ), .A2(\midu/_086_ ), .ZN(\midu/_003_ ) );
OAI21_X1 \midu/_200_ ( .A(\midu/_036_ ), .B1(\midu/_127_ ), .B2(\midu/_085_ ), .ZN(\midu/_087_ ) );
NAND2_X1 \midu/_201_ ( .A1(\midu/_083_ ), .A2(\midu/_087_ ), .ZN(\midu/_004_ ) );
OAI21_X1 \midu/_202_ ( .A(\midu/_037_ ), .B1(\midu/_127_ ), .B2(\midu/_085_ ), .ZN(\midu/_088_ ) );
NAND2_X1 \midu/_203_ ( .A1(\midu/_083_ ), .A2(\midu/_088_ ), .ZN(\midu/_005_ ) );
OAI21_X1 \midu/_204_ ( .A(\midu/_038_ ), .B1(\midu/_127_ ), .B2(\midu/_085_ ), .ZN(\midu/_089_ ) );
NAND2_X1 \midu/_205_ ( .A1(\midu/_083_ ), .A2(\midu/_089_ ), .ZN(\midu/_006_ ) );
OAI21_X1 \midu/_206_ ( .A(\midu/_039_ ), .B1(\midu/_127_ ), .B2(\midu/_085_ ), .ZN(\midu/_090_ ) );
NAND2_X1 \midu/_207_ ( .A1(\midu/_083_ ), .A2(\midu/_090_ ), .ZN(\midu/_007_ ) );
OAI21_X1 \midu/_208_ ( .A(\midu/_040_ ), .B1(\midu/_127_ ), .B2(\midu/_085_ ), .ZN(\midu/_091_ ) );
NAND2_X1 \midu/_209_ ( .A1(\midu/_083_ ), .A2(\midu/_091_ ), .ZN(\midu/_008_ ) );
OAI21_X1 \midu/_210_ ( .A(\midu/_041_ ), .B1(\midu/_127_ ), .B2(\midu/_085_ ), .ZN(\midu/_092_ ) );
NAND2_X1 \midu/_211_ ( .A1(\midu/_083_ ), .A2(\midu/_092_ ), .ZN(\midu/_009_ ) );
OAI21_X1 \midu/_212_ ( .A(\midu/_042_ ), .B1(\midu/_127_ ), .B2(\midu/_085_ ), .ZN(\midu/_093_ ) );
NAND2_X1 \midu/_213_ ( .A1(\midu/_083_ ), .A2(\midu/_093_ ), .ZN(\midu/_010_ ) );
BUF_X4 \midu/_214_ ( .A(\midu/_077_ ), .Z(\midu/_094_ ) );
INV_X1 \midu/_215_ ( .A(\midu/_085_ ), .ZN(\midu/_095_ ) );
BUF_X4 \midu/_216_ ( .A(\midu/_095_ ), .Z(\midu/_096_ ) );
OAI22_X1 \midu/_217_ ( .A1(\midu/_075_ ), .A2(\midu/_094_ ), .B1(\midu/_121_ ), .B2(\midu/_096_ ), .ZN(\midu/_012_ ) );
OAI22_X1 \midu/_218_ ( .A1(\midu/_075_ ), .A2(\midu/_094_ ), .B1(\midu/_130_ ), .B2(\midu/_096_ ), .ZN(\midu/_013_ ) );
OAI22_X1 \midu/_219_ ( .A1(\midu/_075_ ), .A2(\midu/_094_ ), .B1(\midu/_066_ ), .B2(\midu/_096_ ), .ZN(\midu/_014_ ) );
OAI22_X1 \midu/_220_ ( .A1(\midu/_075_ ), .A2(\midu/_094_ ), .B1(\midu/_069_ ), .B2(\midu/_096_ ), .ZN(\midu/_015_ ) );
OAI22_X1 \midu/_221_ ( .A1(\midu/_075_ ), .A2(\midu/_094_ ), .B1(\midu/_072_ ), .B2(\midu/_096_ ), .ZN(\midu/_016_ ) );
OAI22_X1 \midu/_222_ ( .A1(\midu/_075_ ), .A2(\midu/_094_ ), .B1(\midu/_109_ ), .B2(\midu/_096_ ), .ZN(\midu/_017_ ) );
OAI22_X1 \midu/_223_ ( .A1(\midu/_075_ ), .A2(\midu/_094_ ), .B1(\midu/_123_ ), .B2(\midu/_096_ ), .ZN(\midu/_018_ ) );
OAI22_X1 \midu/_224_ ( .A1(\midu/_075_ ), .A2(\midu/_094_ ), .B1(\midu/_065_ ), .B2(\midu/_096_ ), .ZN(\midu/_019_ ) );
OAI22_X1 \midu/_225_ ( .A1(\midu/_074_ ), .A2(\midu/_094_ ), .B1(\midu/_068_ ), .B2(\midu/_096_ ), .ZN(\midu/_020_ ) );
OAI22_X1 \midu/_226_ ( .A1(\midu/_074_ ), .A2(\midu/_094_ ), .B1(\midu/_071_ ), .B2(\midu/_096_ ), .ZN(\midu/_021_ ) );
OAI22_X1 \midu/_227_ ( .A1(\midu/_074_ ), .A2(\midu/_077_ ), .B1(\midu/_076_ ), .B2(\midu/_095_ ), .ZN(\midu/_023_ ) );
AOI21_X1 \midu/_228_ ( .A(\midu/_077_ ), .B1(\midu/_128_ ), .B2(\midu/_095_ ), .ZN(\midu/_097_ ) );
OR3_X2 \midu/_229_ ( .A1(\midu/_081_ ), .A2(\midu/_097_ ), .A3(\midu/_082_ ), .ZN(\midu/_024_ ) );
BUF_X1 \midu/_230_ ( .A(\inst[12] ), .Z(\func[0] ) );
BUF_X1 \midu/_231_ ( .A(\inst[13] ), .Z(\func[1] ) );
BUF_X1 \midu/_232_ ( .A(\inst[14] ), .Z(\func[2] ) );
BUF_X1 \midu/_233_ ( .A(\inst[0] ), .Z(\op[0] ) );
BUF_X1 \midu/_234_ ( .A(\inst[1] ), .Z(\op[1] ) );
BUF_X1 \midu/_235_ ( .A(\inst[2] ), .Z(\op[2] ) );
BUF_X1 \midu/_236_ ( .A(\inst[3] ), .Z(\op[3] ) );
BUF_X1 \midu/_237_ ( .A(\inst[4] ), .Z(\op[4] ) );
BUF_X1 \midu/_238_ ( .A(\inst[5] ), .Z(\op[5] ) );
BUF_X1 \midu/_239_ ( .A(\inst[6] ), .Z(\op[6] ) );
BUF_X1 \midu/_240_ ( .A(\inst[7] ), .Z(\rd[0] ) );
BUF_X1 \midu/_241_ ( .A(\inst[8] ), .Z(\rd[1] ) );
BUF_X1 \midu/_242_ ( .A(\inst[9] ), .Z(\rd[2] ) );
BUF_X1 \midu/_243_ ( .A(\inst[10] ), .Z(\rd[3] ) );
BUF_X1 \midu/_244_ ( .A(\inst[11] ), .Z(\rd[4] ) );
BUF_X1 \midu/_245_ ( .A(\inst[15] ), .Z(\rs1[0] ) );
BUF_X1 \midu/_246_ ( .A(\inst[16] ), .Z(\rs1[1] ) );
BUF_X1 \midu/_247_ ( .A(\inst[17] ), .Z(\rs1[2] ) );
BUF_X1 \midu/_248_ ( .A(\inst[18] ), .Z(\rs1[3] ) );
BUF_X1 \midu/_249_ ( .A(\inst[19] ), .Z(\rs1[4] ) );
BUF_X1 \midu/_250_ ( .A(\inst[20] ), .Z(\rs2[0] ) );
BUF_X1 \midu/_251_ ( .A(\inst[21] ), .Z(\rs2[1] ) );
BUF_X1 \midu/_252_ ( .A(\inst[22] ), .Z(\rs2[2] ) );
BUF_X1 \midu/_253_ ( .A(\inst[23] ), .Z(\rs2[3] ) );
BUF_X1 \midu/_254_ ( .A(\inst[24] ), .Z(\rs2[4] ) );
BUF_X1 \midu/_255_ ( .A(\inst[1] ), .Z(\midu/_043_ ) );
BUF_X1 \midu/_256_ ( .A(\inst[0] ), .Z(\midu/_032_ ) );
BUF_X1 \midu/_257_ ( .A(\inst[3] ), .Z(\midu/_057_ ) );
BUF_X1 \midu/_258_ ( .A(\inst[2] ), .Z(\midu/_054_ ) );
BUF_X1 \midu/_259_ ( .A(\inst[5] ), .Z(\midu/_059_ ) );
BUF_X1 \midu/_260_ ( .A(\inst[4] ), .Z(\midu/_058_ ) );
BUF_X1 \midu/_261_ ( .A(\inst[6] ), .Z(\midu/_060_ ) );
BUF_X1 \midu/_262_ ( .A(\inst[25] ), .Z(\midu/_049_ ) );
BUF_X1 \midu/_263_ ( .A(\inst[7] ), .Z(\midu/_061_ ) );
BUF_X1 \midu/_264_ ( .A(\inst[20] ), .Z(\midu/_044_ ) );
BUF_X1 \midu/_265_ ( .A(\midu/_000_ ), .Z(\imm[0] ) );
BUF_X1 \midu/_266_ ( .A(\inst[26] ), .Z(\midu/_050_ ) );
BUF_X1 \midu/_267_ ( .A(\inst[8] ), .Z(\midu/_062_ ) );
BUF_X1 \midu/_268_ ( .A(\inst[21] ), .Z(\midu/_045_ ) );
BUF_X1 \midu/_269_ ( .A(\midu/_011_ ), .Z(\imm[1] ) );
BUF_X1 \midu/_270_ ( .A(\inst[27] ), .Z(\midu/_051_ ) );
BUF_X1 \midu/_271_ ( .A(\inst[9] ), .Z(\midu/_063_ ) );
BUF_X1 \midu/_272_ ( .A(\inst[22] ), .Z(\midu/_046_ ) );
BUF_X1 \midu/_273_ ( .A(\midu/_022_ ), .Z(\imm[2] ) );
BUF_X1 \midu/_274_ ( .A(\inst[28] ), .Z(\midu/_052_ ) );
BUF_X1 \midu/_275_ ( .A(\inst[10] ), .Z(\midu/_033_ ) );
BUF_X1 \midu/_276_ ( .A(\inst[23] ), .Z(\midu/_047_ ) );
BUF_X1 \midu/_277_ ( .A(\midu/_025_ ), .Z(\imm[3] ) );
BUF_X1 \midu/_278_ ( .A(\inst[29] ), .Z(\midu/_053_ ) );
BUF_X1 \midu/_279_ ( .A(\inst[11] ), .Z(\midu/_034_ ) );
BUF_X1 \midu/_280_ ( .A(\inst[24] ), .Z(\midu/_048_ ) );
BUF_X1 \midu/_281_ ( .A(\midu/_026_ ), .Z(\imm[4] ) );
BUF_X1 \midu/_282_ ( .A(\inst[30] ), .Z(\midu/_055_ ) );
BUF_X1 \midu/_283_ ( .A(\midu/_027_ ), .Z(\imm[5] ) );
BUF_X1 \midu/_284_ ( .A(\inst[31] ), .Z(\midu/_056_ ) );
BUF_X1 \midu/_285_ ( .A(\midu/_028_ ), .Z(\imm[6] ) );
BUF_X1 \midu/_286_ ( .A(\midu/_029_ ), .Z(\imm[7] ) );
BUF_X1 \midu/_287_ ( .A(\midu/_030_ ), .Z(\imm[8] ) );
BUF_X1 \midu/_288_ ( .A(\midu/_031_ ), .Z(\imm[9] ) );
BUF_X1 \midu/_289_ ( .A(\midu/_001_ ), .Z(\imm[10] ) );
BUF_X1 \midu/_290_ ( .A(\midu/_002_ ), .Z(\imm[11] ) );
BUF_X1 \midu/_291_ ( .A(\inst[12] ), .Z(\midu/_035_ ) );
BUF_X1 \midu/_292_ ( .A(\midu/_003_ ), .Z(\imm[12] ) );
BUF_X1 \midu/_293_ ( .A(\inst[13] ), .Z(\midu/_036_ ) );
BUF_X1 \midu/_294_ ( .A(\midu/_004_ ), .Z(\imm[13] ) );
BUF_X1 \midu/_295_ ( .A(\inst[14] ), .Z(\midu/_037_ ) );
BUF_X1 \midu/_296_ ( .A(\midu/_005_ ), .Z(\imm[14] ) );
BUF_X1 \midu/_297_ ( .A(\inst[15] ), .Z(\midu/_038_ ) );
BUF_X1 \midu/_298_ ( .A(\midu/_006_ ), .Z(\imm[15] ) );
BUF_X1 \midu/_299_ ( .A(\inst[16] ), .Z(\midu/_039_ ) );
BUF_X1 \midu/_300_ ( .A(\midu/_007_ ), .Z(\imm[16] ) );
BUF_X1 \midu/_301_ ( .A(\inst[17] ), .Z(\midu/_040_ ) );
BUF_X1 \midu/_302_ ( .A(\midu/_008_ ), .Z(\imm[17] ) );
BUF_X1 \midu/_303_ ( .A(\inst[18] ), .Z(\midu/_041_ ) );
BUF_X1 \midu/_304_ ( .A(\midu/_009_ ), .Z(\imm[18] ) );
BUF_X1 \midu/_305_ ( .A(\inst[19] ), .Z(\midu/_042_ ) );
BUF_X1 \midu/_306_ ( .A(\midu/_010_ ), .Z(\imm[19] ) );
BUF_X1 \midu/_307_ ( .A(\midu/_012_ ), .Z(\imm[20] ) );
BUF_X1 \midu/_308_ ( .A(\midu/_013_ ), .Z(\imm[21] ) );
BUF_X1 \midu/_309_ ( .A(\midu/_014_ ), .Z(\imm[22] ) );
BUF_X1 \midu/_310_ ( .A(\midu/_015_ ), .Z(\imm[23] ) );
BUF_X1 \midu/_311_ ( .A(\midu/_016_ ), .Z(\imm[24] ) );
BUF_X1 \midu/_312_ ( .A(\midu/_017_ ), .Z(\imm[25] ) );
BUF_X1 \midu/_313_ ( .A(\midu/_018_ ), .Z(\imm[26] ) );
BUF_X1 \midu/_314_ ( .A(\midu/_019_ ), .Z(\imm[27] ) );
BUF_X1 \midu/_315_ ( .A(\midu/_020_ ), .Z(\imm[28] ) );
BUF_X1 \midu/_316_ ( .A(\midu/_021_ ), .Z(\imm[29] ) );
BUF_X1 \midu/_317_ ( .A(\midu/_023_ ), .Z(\imm[30] ) );
BUF_X1 \midu/_318_ ( .A(\midu/_024_ ), .Z(\imm[31] ) );
INV_X1 \mifu/_224_ ( .A(\mifu/_151_ ), .ZN(\mifu/_106_ ) );
CLKBUF_X2 \mifu/_225_ ( .A(\mifu/_106_ ), .Z(\mifu/_107_ ) );
AND2_X1 \mifu/_226_ ( .A1(\mifu/_107_ ), .A2(\mifu/_072_ ), .ZN(\mifu/_002_ ) );
INV_X1 \mifu/_227_ ( .A(\mifu/_152_ ), .ZN(\mifu/_108_ ) );
NOR3_X1 \mifu/_228_ ( .A1(\mifu/_108_ ), .A2(\mifu/_039_ ), .A3(\mifu/_105_ ), .ZN(\mifu/_109_ ) );
OR3_X4 \mifu/_229_ ( .A1(\mifu/_108_ ), .A2(\mifu/_038_ ), .A3(\mifu/_105_ ), .ZN(\mifu/_110_ ) );
INV_X1 \mifu/_230_ ( .A(\mifu/_001_ ), .ZN(\mifu/_111_ ) );
AOI211_X2 \mifu/_231_ ( .A(\mifu/_151_ ), .B(\mifu/_109_ ), .C1(\mifu/_110_ ), .C2(\mifu/_111_ ), .ZN(\mifu/_003_ ) );
AND2_X4 \mifu/_232_ ( .A1(\mifu/_039_ ), .A2(\mifu/_038_ ), .ZN(\mifu/_112_ ) );
MUX2_X1 \mifu/_233_ ( .A(\mifu/_105_ ), .B(\mifu/_150_ ), .S(\mifu/_112_ ), .Z(\mifu/_113_ ) );
AND3_X1 \mifu/_234_ ( .A1(\mifu/_113_ ), .A2(\mifu/_106_ ), .A3(\mifu/_152_ ), .ZN(\mifu/_004_ ) );
MUX2_X1 \mifu/_235_ ( .A(\mifu/_073_ ), .B(\mifu/_040_ ), .S(\mifu/_072_ ), .Z(\mifu/_114_ ) );
AND2_X1 \mifu/_236_ ( .A1(\mifu/_114_ ), .A2(\mifu/_107_ ), .ZN(\mifu/_005_ ) );
MUX2_X1 \mifu/_237_ ( .A(\mifu/_084_ ), .B(\mifu/_051_ ), .S(\mifu/_072_ ), .Z(\mifu/_115_ ) );
AND2_X1 \mifu/_238_ ( .A1(\mifu/_115_ ), .A2(\mifu/_107_ ), .ZN(\mifu/_006_ ) );
MUX2_X1 \mifu/_239_ ( .A(\mifu/_095_ ), .B(\mifu/_062_ ), .S(\mifu/_072_ ), .Z(\mifu/_116_ ) );
AND2_X1 \mifu/_240_ ( .A1(\mifu/_116_ ), .A2(\mifu/_107_ ), .ZN(\mifu/_007_ ) );
MUX2_X1 \mifu/_241_ ( .A(\mifu/_098_ ), .B(\mifu/_065_ ), .S(\mifu/_072_ ), .Z(\mifu/_117_ ) );
AND2_X1 \mifu/_242_ ( .A1(\mifu/_117_ ), .A2(\mifu/_107_ ), .ZN(\mifu/_008_ ) );
MUX2_X1 \mifu/_243_ ( .A(\mifu/_099_ ), .B(\mifu/_066_ ), .S(\mifu/_072_ ), .Z(\mifu/_118_ ) );
AND2_X1 \mifu/_244_ ( .A1(\mifu/_118_ ), .A2(\mifu/_107_ ), .ZN(\mifu/_009_ ) );
MUX2_X1 \mifu/_245_ ( .A(\mifu/_100_ ), .B(\mifu/_067_ ), .S(\mifu/_072_ ), .Z(\mifu/_119_ ) );
AND2_X1 \mifu/_246_ ( .A1(\mifu/_119_ ), .A2(\mifu/_107_ ), .ZN(\mifu/_010_ ) );
MUX2_X1 \mifu/_247_ ( .A(\mifu/_101_ ), .B(\mifu/_068_ ), .S(\mifu/_072_ ), .Z(\mifu/_120_ ) );
AND2_X1 \mifu/_248_ ( .A1(\mifu/_120_ ), .A2(\mifu/_107_ ), .ZN(\mifu/_011_ ) );
MUX2_X1 \mifu/_249_ ( .A(\mifu/_102_ ), .B(\mifu/_069_ ), .S(\mifu/_072_ ), .Z(\mifu/_121_ ) );
AND2_X1 \mifu/_250_ ( .A1(\mifu/_121_ ), .A2(\mifu/_107_ ), .ZN(\mifu/_012_ ) );
MUX2_X1 \mifu/_251_ ( .A(\mifu/_103_ ), .B(\mifu/_070_ ), .S(\mifu/_072_ ), .Z(\mifu/_122_ ) );
AND2_X1 \mifu/_252_ ( .A1(\mifu/_122_ ), .A2(\mifu/_107_ ), .ZN(\mifu/_013_ ) );
MUX2_X1 \mifu/_253_ ( .A(\mifu/_104_ ), .B(\mifu/_071_ ), .S(\mifu/_072_ ), .Z(\mifu/_123_ ) );
CLKBUF_X2 \mifu/_254_ ( .A(\mifu/_106_ ), .Z(\mifu/_124_ ) );
AND2_X1 \mifu/_255_ ( .A1(\mifu/_123_ ), .A2(\mifu/_124_ ), .ZN(\mifu/_014_ ) );
MUX2_X1 \mifu/_256_ ( .A(\mifu/_074_ ), .B(\mifu/_041_ ), .S(\mifu/_072_ ), .Z(\mifu/_125_ ) );
AND2_X1 \mifu/_257_ ( .A1(\mifu/_125_ ), .A2(\mifu/_124_ ), .ZN(\mifu/_015_ ) );
MUX2_X1 \mifu/_258_ ( .A(\mifu/_075_ ), .B(\mifu/_042_ ), .S(\mifu/_072_ ), .Z(\mifu/_126_ ) );
AND2_X1 \mifu/_259_ ( .A1(\mifu/_126_ ), .A2(\mifu/_124_ ), .ZN(\mifu/_016_ ) );
MUX2_X1 \mifu/_260_ ( .A(\mifu/_076_ ), .B(\mifu/_043_ ), .S(\mifu/_072_ ), .Z(\mifu/_127_ ) );
AND2_X1 \mifu/_261_ ( .A1(\mifu/_127_ ), .A2(\mifu/_124_ ), .ZN(\mifu/_017_ ) );
MUX2_X1 \mifu/_262_ ( .A(\mifu/_077_ ), .B(\mifu/_044_ ), .S(\mifu/_072_ ), .Z(\mifu/_128_ ) );
AND2_X1 \mifu/_263_ ( .A1(\mifu/_128_ ), .A2(\mifu/_124_ ), .ZN(\mifu/_018_ ) );
MUX2_X1 \mifu/_264_ ( .A(\mifu/_078_ ), .B(\mifu/_045_ ), .S(\mifu/_072_ ), .Z(\mifu/_129_ ) );
AND2_X1 \mifu/_265_ ( .A1(\mifu/_129_ ), .A2(\mifu/_124_ ), .ZN(\mifu/_019_ ) );
MUX2_X1 \mifu/_266_ ( .A(\mifu/_079_ ), .B(\mifu/_046_ ), .S(\mifu/_072_ ), .Z(\mifu/_130_ ) );
AND2_X1 \mifu/_267_ ( .A1(\mifu/_130_ ), .A2(\mifu/_124_ ), .ZN(\mifu/_020_ ) );
MUX2_X1 \mifu/_268_ ( .A(\mifu/_080_ ), .B(\mifu/_047_ ), .S(\mifu/_072_ ), .Z(\mifu/_131_ ) );
AND2_X1 \mifu/_269_ ( .A1(\mifu/_131_ ), .A2(\mifu/_124_ ), .ZN(\mifu/_021_ ) );
MUX2_X1 \mifu/_270_ ( .A(\mifu/_081_ ), .B(\mifu/_048_ ), .S(\mifu/_072_ ), .Z(\mifu/_132_ ) );
AND2_X1 \mifu/_271_ ( .A1(\mifu/_132_ ), .A2(\mifu/_124_ ), .ZN(\mifu/_022_ ) );
MUX2_X1 \mifu/_272_ ( .A(\mifu/_082_ ), .B(\mifu/_049_ ), .S(\mifu/_072_ ), .Z(\mifu/_133_ ) );
AND2_X1 \mifu/_273_ ( .A1(\mifu/_133_ ), .A2(\mifu/_124_ ), .ZN(\mifu/_023_ ) );
MUX2_X1 \mifu/_274_ ( .A(\mifu/_083_ ), .B(\mifu/_050_ ), .S(\mifu/_072_ ), .Z(\mifu/_134_ ) );
CLKBUF_X2 \mifu/_275_ ( .A(\mifu/_106_ ), .Z(\mifu/_135_ ) );
AND2_X1 \mifu/_276_ ( .A1(\mifu/_134_ ), .A2(\mifu/_135_ ), .ZN(\mifu/_024_ ) );
MUX2_X1 \mifu/_277_ ( .A(\mifu/_085_ ), .B(\mifu/_052_ ), .S(\mifu/_072_ ), .Z(\mifu/_136_ ) );
AND2_X1 \mifu/_278_ ( .A1(\mifu/_136_ ), .A2(\mifu/_135_ ), .ZN(\mifu/_025_ ) );
MUX2_X1 \mifu/_279_ ( .A(\mifu/_086_ ), .B(\mifu/_053_ ), .S(\mifu/_072_ ), .Z(\mifu/_137_ ) );
AND2_X1 \mifu/_280_ ( .A1(\mifu/_137_ ), .A2(\mifu/_135_ ), .ZN(\mifu/_026_ ) );
MUX2_X1 \mifu/_281_ ( .A(\mifu/_087_ ), .B(\mifu/_054_ ), .S(\mifu/_072_ ), .Z(\mifu/_138_ ) );
AND2_X1 \mifu/_282_ ( .A1(\mifu/_138_ ), .A2(\mifu/_135_ ), .ZN(\mifu/_027_ ) );
MUX2_X1 \mifu/_283_ ( .A(\mifu/_088_ ), .B(\mifu/_055_ ), .S(\mifu/_072_ ), .Z(\mifu/_139_ ) );
AND2_X1 \mifu/_284_ ( .A1(\mifu/_139_ ), .A2(\mifu/_135_ ), .ZN(\mifu/_028_ ) );
MUX2_X1 \mifu/_285_ ( .A(\mifu/_089_ ), .B(\mifu/_056_ ), .S(\mifu/_072_ ), .Z(\mifu/_140_ ) );
AND2_X1 \mifu/_286_ ( .A1(\mifu/_140_ ), .A2(\mifu/_135_ ), .ZN(\mifu/_029_ ) );
MUX2_X1 \mifu/_287_ ( .A(\mifu/_090_ ), .B(\mifu/_057_ ), .S(\mifu/_072_ ), .Z(\mifu/_141_ ) );
AND2_X1 \mifu/_288_ ( .A1(\mifu/_141_ ), .A2(\mifu/_135_ ), .ZN(\mifu/_030_ ) );
MUX2_X1 \mifu/_289_ ( .A(\mifu/_091_ ), .B(\mifu/_058_ ), .S(\mifu/_072_ ), .Z(\mifu/_142_ ) );
AND2_X1 \mifu/_290_ ( .A1(\mifu/_142_ ), .A2(\mifu/_135_ ), .ZN(\mifu/_031_ ) );
MUX2_X1 \mifu/_291_ ( .A(\mifu/_092_ ), .B(\mifu/_059_ ), .S(\mifu/_072_ ), .Z(\mifu/_143_ ) );
AND2_X1 \mifu/_292_ ( .A1(\mifu/_143_ ), .A2(\mifu/_135_ ), .ZN(\mifu/_032_ ) );
MUX2_X1 \mifu/_293_ ( .A(\mifu/_093_ ), .B(\mifu/_060_ ), .S(\mifu/_072_ ), .Z(\mifu/_144_ ) );
AND2_X1 \mifu/_294_ ( .A1(\mifu/_144_ ), .A2(\mifu/_135_ ), .ZN(\mifu/_033_ ) );
MUX2_X1 \mifu/_295_ ( .A(\mifu/_094_ ), .B(\mifu/_061_ ), .S(\mifu/_072_ ), .Z(\mifu/_145_ ) );
AND2_X1 \mifu/_296_ ( .A1(\mifu/_145_ ), .A2(\mifu/_106_ ), .ZN(\mifu/_034_ ) );
MUX2_X1 \mifu/_297_ ( .A(\mifu/_096_ ), .B(\mifu/_063_ ), .S(\mifu/_072_ ), .Z(\mifu/_146_ ) );
AND2_X1 \mifu/_298_ ( .A1(\mifu/_146_ ), .A2(\mifu/_106_ ), .ZN(\mifu/_035_ ) );
MUX2_X1 \mifu/_299_ ( .A(\mifu/_097_ ), .B(\mifu/_064_ ), .S(\mifu/_072_ ), .Z(\mifu/_147_ ) );
AND2_X1 \mifu/_300_ ( .A1(\mifu/_147_ ), .A2(\mifu/_106_ ), .ZN(\mifu/_036_ ) );
INV_X1 \mifu/_301_ ( .A(\mifu/_112_ ), .ZN(\mifu/_148_ ) );
NAND3_X1 \mifu/_302_ ( .A1(\mifu/_148_ ), .A2(\mifu/_105_ ), .A3(\mifu/_111_ ), .ZN(\mifu/_149_ ) );
AND2_X1 \mifu/_303_ ( .A1(\mifu/_149_ ), .A2(\mifu/_106_ ), .ZN(\mifu/_037_ ) );
DFF_X1 \mifu/_304_ ( .CK(clk ), .D(\mifu/_188_ ), .Q(inst_valid ), .QN(\mifu/_187_ ) );
DFF_X1 \mifu/_305_ ( .CK(clk ), .D(\mifu/_189_ ), .Q(ifu_arvalid ), .QN(\mifu/_186_ ) );
DFF_X1 \mifu/_306_ ( .CK(clk ), .D(\mifu/_190_ ), .Q(pc_wen ), .QN(\mifu/_185_ ) );
DFF_X1 \mifu/_307_ ( .CK(clk ), .D(\mifu/_191_ ), .Q(\inst[0] ), .QN(\mifu/_184_ ) );
DFF_X1 \mifu/_308_ ( .CK(clk ), .D(\mifu/_192_ ), .Q(\inst[1] ), .QN(\mifu/_183_ ) );
DFF_X1 \mifu/_309_ ( .CK(clk ), .D(\mifu/_193_ ), .Q(\inst[2] ), .QN(\mifu/_182_ ) );
DFF_X1 \mifu/_310_ ( .CK(clk ), .D(\mifu/_194_ ), .Q(\inst[3] ), .QN(\mifu/_181_ ) );
DFF_X1 \mifu/_311_ ( .CK(clk ), .D(\mifu/_195_ ), .Q(\inst[4] ), .QN(\mifu/_180_ ) );
DFF_X1 \mifu/_312_ ( .CK(clk ), .D(\mifu/_196_ ), .Q(\inst[5] ), .QN(\mifu/_179_ ) );
DFF_X1 \mifu/_313_ ( .CK(clk ), .D(\mifu/_197_ ), .Q(\inst[6] ), .QN(\mifu/_178_ ) );
DFF_X1 \mifu/_314_ ( .CK(clk ), .D(\mifu/_198_ ), .Q(\inst[7] ), .QN(\mifu/_177_ ) );
DFF_X1 \mifu/_315_ ( .CK(clk ), .D(\mifu/_199_ ), .Q(\inst[8] ), .QN(\mifu/_176_ ) );
DFF_X1 \mifu/_316_ ( .CK(clk ), .D(\mifu/_200_ ), .Q(\inst[9] ), .QN(\mifu/_175_ ) );
DFF_X1 \mifu/_317_ ( .CK(clk ), .D(\mifu/_201_ ), .Q(\inst[10] ), .QN(\mifu/_174_ ) );
DFF_X1 \mifu/_318_ ( .CK(clk ), .D(\mifu/_202_ ), .Q(\inst[11] ), .QN(\mifu/_173_ ) );
DFF_X1 \mifu/_319_ ( .CK(clk ), .D(\mifu/_203_ ), .Q(\inst[12] ), .QN(\mifu/_172_ ) );
DFF_X1 \mifu/_320_ ( .CK(clk ), .D(\mifu/_204_ ), .Q(\inst[13] ), .QN(\mifu/_171_ ) );
DFF_X1 \mifu/_321_ ( .CK(clk ), .D(\mifu/_205_ ), .Q(\inst[14] ), .QN(\mifu/_170_ ) );
DFF_X1 \mifu/_322_ ( .CK(clk ), .D(\mifu/_206_ ), .Q(\inst[15] ), .QN(\mifu/_169_ ) );
DFF_X1 \mifu/_323_ ( .CK(clk ), .D(\mifu/_207_ ), .Q(\inst[16] ), .QN(\mifu/_168_ ) );
DFF_X1 \mifu/_324_ ( .CK(clk ), .D(\mifu/_208_ ), .Q(\inst[17] ), .QN(\mifu/_167_ ) );
DFF_X1 \mifu/_325_ ( .CK(clk ), .D(\mifu/_209_ ), .Q(\inst[18] ), .QN(\mifu/_166_ ) );
DFF_X1 \mifu/_326_ ( .CK(clk ), .D(\mifu/_210_ ), .Q(\inst[19] ), .QN(\mifu/_165_ ) );
DFF_X1 \mifu/_327_ ( .CK(clk ), .D(\mifu/_211_ ), .Q(\inst[20] ), .QN(\mifu/_164_ ) );
DFF_X1 \mifu/_328_ ( .CK(clk ), .D(\mifu/_212_ ), .Q(\inst[21] ), .QN(\mifu/_163_ ) );
DFF_X1 \mifu/_329_ ( .CK(clk ), .D(\mifu/_213_ ), .Q(\inst[22] ), .QN(\mifu/_162_ ) );
DFF_X1 \mifu/_330_ ( .CK(clk ), .D(\mifu/_214_ ), .Q(\inst[23] ), .QN(\mifu/_161_ ) );
DFF_X1 \mifu/_331_ ( .CK(clk ), .D(\mifu/_215_ ), .Q(\inst[24] ), .QN(\mifu/_160_ ) );
DFF_X1 \mifu/_332_ ( .CK(clk ), .D(\mifu/_216_ ), .Q(\inst[25] ), .QN(\mifu/_159_ ) );
DFF_X1 \mifu/_333_ ( .CK(clk ), .D(\mifu/_217_ ), .Q(\inst[26] ), .QN(\mifu/_158_ ) );
DFF_X1 \mifu/_334_ ( .CK(clk ), .D(\mifu/_218_ ), .Q(\inst[27] ), .QN(\mifu/_157_ ) );
DFF_X1 \mifu/_335_ ( .CK(clk ), .D(\mifu/_219_ ), .Q(\inst[28] ), .QN(\mifu/_156_ ) );
DFF_X1 \mifu/_336_ ( .CK(clk ), .D(\mifu/_220_ ), .Q(\inst[29] ), .QN(\mifu/_155_ ) );
DFF_X1 \mifu/_337_ ( .CK(clk ), .D(\mifu/_221_ ), .Q(\inst[30] ), .QN(\mifu/_154_ ) );
DFF_X1 \mifu/_338_ ( .CK(clk ), .D(\mifu/_222_ ), .Q(\inst[31] ), .QN(\mifu/_153_ ) );
DFF_X1 \mifu/_339_ ( .CK(clk ), .D(\mifu/_223_ ), .Q(\mifu/wait_ready ), .QN(\mifu/_000_ ) );
BUF_X1 \mifu/_340_ ( .A(\pc[0] ), .Z(\ifu_araddr[0] ) );
BUF_X1 \mifu/_341_ ( .A(\pc[1] ), .Z(\ifu_araddr[1] ) );
BUF_X1 \mifu/_342_ ( .A(\pc[2] ), .Z(\ifu_araddr[2] ) );
BUF_X1 \mifu/_343_ ( .A(\pc[3] ), .Z(\ifu_araddr[3] ) );
BUF_X1 \mifu/_344_ ( .A(\pc[4] ), .Z(\ifu_araddr[4] ) );
BUF_X1 \mifu/_345_ ( .A(\pc[5] ), .Z(\ifu_araddr[5] ) );
BUF_X1 \mifu/_346_ ( .A(\pc[6] ), .Z(\ifu_araddr[6] ) );
BUF_X1 \mifu/_347_ ( .A(\pc[7] ), .Z(\ifu_araddr[7] ) );
BUF_X1 \mifu/_348_ ( .A(\pc[8] ), .Z(\ifu_araddr[8] ) );
BUF_X1 \mifu/_349_ ( .A(\pc[9] ), .Z(\ifu_araddr[9] ) );
BUF_X1 \mifu/_350_ ( .A(\pc[10] ), .Z(\ifu_araddr[10] ) );
BUF_X1 \mifu/_351_ ( .A(\pc[11] ), .Z(\ifu_araddr[11] ) );
BUF_X1 \mifu/_352_ ( .A(\pc[12] ), .Z(\ifu_araddr[12] ) );
BUF_X1 \mifu/_353_ ( .A(\pc[13] ), .Z(\ifu_araddr[13] ) );
BUF_X1 \mifu/_354_ ( .A(\pc[14] ), .Z(\ifu_araddr[14] ) );
BUF_X1 \mifu/_355_ ( .A(\pc[15] ), .Z(\ifu_araddr[15] ) );
BUF_X1 \mifu/_356_ ( .A(\pc[16] ), .Z(\ifu_araddr[16] ) );
BUF_X1 \mifu/_357_ ( .A(\pc[17] ), .Z(\ifu_araddr[17] ) );
BUF_X1 \mifu/_358_ ( .A(\pc[18] ), .Z(\ifu_araddr[18] ) );
BUF_X1 \mifu/_359_ ( .A(\pc[19] ), .Z(\ifu_araddr[19] ) );
BUF_X1 \mifu/_360_ ( .A(\pc[20] ), .Z(\ifu_araddr[20] ) );
BUF_X1 \mifu/_361_ ( .A(\pc[21] ), .Z(\ifu_araddr[21] ) );
BUF_X1 \mifu/_362_ ( .A(\pc[22] ), .Z(\ifu_araddr[22] ) );
BUF_X1 \mifu/_363_ ( .A(\pc[23] ), .Z(\ifu_araddr[23] ) );
BUF_X1 \mifu/_364_ ( .A(\pc[24] ), .Z(\ifu_araddr[24] ) );
BUF_X1 \mifu/_365_ ( .A(\pc[25] ), .Z(\ifu_araddr[25] ) );
BUF_X1 \mifu/_366_ ( .A(\pc[26] ), .Z(\ifu_araddr[26] ) );
BUF_X1 \mifu/_367_ ( .A(\pc[27] ), .Z(\ifu_araddr[27] ) );
BUF_X1 \mifu/_368_ ( .A(\pc[28] ), .Z(\ifu_araddr[28] ) );
BUF_X1 \mifu/_369_ ( .A(\pc[29] ), .Z(\ifu_araddr[29] ) );
BUF_X1 \mifu/_370_ ( .A(\pc[30] ), .Z(\ifu_araddr[30] ) );
BUF_X1 \mifu/_371_ ( .A(\pc[31] ), .Z(\ifu_araddr[31] ) );
BUF_X1 \mifu/_372_ ( .A(1'b0 ), .Z(ifu_rready ) );
BUF_X1 \mifu/_373_ ( .A(rst ), .Z(\mifu/_151_ ) );
BUF_X1 \mifu/_374_ ( .A(\mifu/wait_ready ), .Z(\mifu/_152_ ) );
BUF_X1 \mifu/_375_ ( .A(ifu_arvalid ), .Z(\mifu/_039_ ) );
BUF_X1 \mifu/_376_ ( .A(ifu_arready ), .Z(\mifu/_038_ ) );
BUF_X1 \mifu/_377_ ( .A(lsu_finish ), .Z(\mifu/_105_ ) );
BUF_X1 \mifu/_378_ ( .A(\mifu/_000_ ), .Z(\mifu/_001_ ) );
BUF_X1 \mifu/_379_ ( .A(\inst[0] ), .Z(\mifu/_073_ ) );
BUF_X1 \mifu/_380_ ( .A(\ifu_rdata[0] ), .Z(\mifu/_040_ ) );
BUF_X1 \mifu/_381_ ( .A(ifu_rvalid ), .Z(\mifu/_072_ ) );
BUF_X1 \mifu/_382_ ( .A(\inst[1] ), .Z(\mifu/_084_ ) );
BUF_X1 \mifu/_383_ ( .A(\ifu_rdata[1] ), .Z(\mifu/_051_ ) );
BUF_X1 \mifu/_384_ ( .A(\inst[2] ), .Z(\mifu/_095_ ) );
BUF_X1 \mifu/_385_ ( .A(\ifu_rdata[2] ), .Z(\mifu/_062_ ) );
BUF_X1 \mifu/_386_ ( .A(\inst[3] ), .Z(\mifu/_098_ ) );
BUF_X1 \mifu/_387_ ( .A(\ifu_rdata[3] ), .Z(\mifu/_065_ ) );
BUF_X1 \mifu/_388_ ( .A(\inst[4] ), .Z(\mifu/_099_ ) );
BUF_X1 \mifu/_389_ ( .A(\ifu_rdata[4] ), .Z(\mifu/_066_ ) );
BUF_X1 \mifu/_390_ ( .A(\inst[5] ), .Z(\mifu/_100_ ) );
BUF_X1 \mifu/_391_ ( .A(\ifu_rdata[5] ), .Z(\mifu/_067_ ) );
BUF_X1 \mifu/_392_ ( .A(\inst[6] ), .Z(\mifu/_101_ ) );
BUF_X1 \mifu/_393_ ( .A(\ifu_rdata[6] ), .Z(\mifu/_068_ ) );
BUF_X1 \mifu/_394_ ( .A(\inst[7] ), .Z(\mifu/_102_ ) );
BUF_X1 \mifu/_395_ ( .A(\ifu_rdata[7] ), .Z(\mifu/_069_ ) );
BUF_X1 \mifu/_396_ ( .A(\inst[8] ), .Z(\mifu/_103_ ) );
BUF_X1 \mifu/_397_ ( .A(\ifu_rdata[8] ), .Z(\mifu/_070_ ) );
BUF_X1 \mifu/_398_ ( .A(\inst[9] ), .Z(\mifu/_104_ ) );
BUF_X1 \mifu/_399_ ( .A(\ifu_rdata[9] ), .Z(\mifu/_071_ ) );
BUF_X1 \mifu/_400_ ( .A(\inst[10] ), .Z(\mifu/_074_ ) );
BUF_X1 \mifu/_401_ ( .A(\ifu_rdata[10] ), .Z(\mifu/_041_ ) );
BUF_X1 \mifu/_402_ ( .A(\inst[11] ), .Z(\mifu/_075_ ) );
BUF_X1 \mifu/_403_ ( .A(\ifu_rdata[11] ), .Z(\mifu/_042_ ) );
BUF_X1 \mifu/_404_ ( .A(\inst[12] ), .Z(\mifu/_076_ ) );
BUF_X1 \mifu/_405_ ( .A(\ifu_rdata[12] ), .Z(\mifu/_043_ ) );
BUF_X1 \mifu/_406_ ( .A(\inst[13] ), .Z(\mifu/_077_ ) );
BUF_X1 \mifu/_407_ ( .A(\ifu_rdata[13] ), .Z(\mifu/_044_ ) );
BUF_X1 \mifu/_408_ ( .A(\inst[14] ), .Z(\mifu/_078_ ) );
BUF_X1 \mifu/_409_ ( .A(\ifu_rdata[14] ), .Z(\mifu/_045_ ) );
BUF_X1 \mifu/_410_ ( .A(\inst[15] ), .Z(\mifu/_079_ ) );
BUF_X1 \mifu/_411_ ( .A(\ifu_rdata[15] ), .Z(\mifu/_046_ ) );
BUF_X1 \mifu/_412_ ( .A(\inst[16] ), .Z(\mifu/_080_ ) );
BUF_X1 \mifu/_413_ ( .A(\ifu_rdata[16] ), .Z(\mifu/_047_ ) );
BUF_X1 \mifu/_414_ ( .A(\inst[17] ), .Z(\mifu/_081_ ) );
BUF_X1 \mifu/_415_ ( .A(\ifu_rdata[17] ), .Z(\mifu/_048_ ) );
BUF_X1 \mifu/_416_ ( .A(\inst[18] ), .Z(\mifu/_082_ ) );
BUF_X1 \mifu/_417_ ( .A(\ifu_rdata[18] ), .Z(\mifu/_049_ ) );
BUF_X1 \mifu/_418_ ( .A(\inst[19] ), .Z(\mifu/_083_ ) );
BUF_X1 \mifu/_419_ ( .A(\ifu_rdata[19] ), .Z(\mifu/_050_ ) );
BUF_X1 \mifu/_420_ ( .A(\inst[20] ), .Z(\mifu/_085_ ) );
BUF_X1 \mifu/_421_ ( .A(\ifu_rdata[20] ), .Z(\mifu/_052_ ) );
BUF_X1 \mifu/_422_ ( .A(\inst[21] ), .Z(\mifu/_086_ ) );
BUF_X1 \mifu/_423_ ( .A(\ifu_rdata[21] ), .Z(\mifu/_053_ ) );
BUF_X1 \mifu/_424_ ( .A(\inst[22] ), .Z(\mifu/_087_ ) );
BUF_X1 \mifu/_425_ ( .A(\ifu_rdata[22] ), .Z(\mifu/_054_ ) );
BUF_X1 \mifu/_426_ ( .A(\inst[23] ), .Z(\mifu/_088_ ) );
BUF_X1 \mifu/_427_ ( .A(\ifu_rdata[23] ), .Z(\mifu/_055_ ) );
BUF_X1 \mifu/_428_ ( .A(\inst[24] ), .Z(\mifu/_089_ ) );
BUF_X1 \mifu/_429_ ( .A(\ifu_rdata[24] ), .Z(\mifu/_056_ ) );
BUF_X1 \mifu/_430_ ( .A(\inst[25] ), .Z(\mifu/_090_ ) );
BUF_X1 \mifu/_431_ ( .A(\ifu_rdata[25] ), .Z(\mifu/_057_ ) );
BUF_X1 \mifu/_432_ ( .A(\inst[26] ), .Z(\mifu/_091_ ) );
BUF_X1 \mifu/_433_ ( .A(\ifu_rdata[26] ), .Z(\mifu/_058_ ) );
BUF_X1 \mifu/_434_ ( .A(\inst[27] ), .Z(\mifu/_092_ ) );
BUF_X1 \mifu/_435_ ( .A(\ifu_rdata[27] ), .Z(\mifu/_059_ ) );
BUF_X1 \mifu/_436_ ( .A(\inst[28] ), .Z(\mifu/_093_ ) );
BUF_X1 \mifu/_437_ ( .A(\ifu_rdata[28] ), .Z(\mifu/_060_ ) );
BUF_X1 \mifu/_438_ ( .A(\inst[29] ), .Z(\mifu/_094_ ) );
BUF_X1 \mifu/_439_ ( .A(\ifu_rdata[29] ), .Z(\mifu/_061_ ) );
BUF_X1 \mifu/_440_ ( .A(\inst[30] ), .Z(\mifu/_096_ ) );
BUF_X1 \mifu/_441_ ( .A(\ifu_rdata[30] ), .Z(\mifu/_063_ ) );
BUF_X1 \mifu/_442_ ( .A(\inst[31] ), .Z(\mifu/_097_ ) );
BUF_X1 \mifu/_443_ ( .A(\ifu_rdata[31] ), .Z(\mifu/_064_ ) );
BUF_X1 \mifu/_444_ ( .A(pc_wen ), .Z(\mifu/_150_ ) );
BUF_X1 \mifu/_445_ ( .A(\mifu/_002_ ), .Z(\mifu/_188_ ) );
BUF_X1 \mifu/_446_ ( .A(\mifu/_003_ ), .Z(\mifu/_189_ ) );
BUF_X1 \mifu/_447_ ( .A(\mifu/_004_ ), .Z(\mifu/_190_ ) );
BUF_X1 \mifu/_448_ ( .A(\mifu/_005_ ), .Z(\mifu/_191_ ) );
BUF_X1 \mifu/_449_ ( .A(\mifu/_006_ ), .Z(\mifu/_192_ ) );
BUF_X1 \mifu/_450_ ( .A(\mifu/_007_ ), .Z(\mifu/_193_ ) );
BUF_X1 \mifu/_451_ ( .A(\mifu/_008_ ), .Z(\mifu/_194_ ) );
BUF_X1 \mifu/_452_ ( .A(\mifu/_009_ ), .Z(\mifu/_195_ ) );
BUF_X1 \mifu/_453_ ( .A(\mifu/_010_ ), .Z(\mifu/_196_ ) );
BUF_X1 \mifu/_454_ ( .A(\mifu/_011_ ), .Z(\mifu/_197_ ) );
BUF_X1 \mifu/_455_ ( .A(\mifu/_012_ ), .Z(\mifu/_198_ ) );
BUF_X1 \mifu/_456_ ( .A(\mifu/_013_ ), .Z(\mifu/_199_ ) );
BUF_X1 \mifu/_457_ ( .A(\mifu/_014_ ), .Z(\mifu/_200_ ) );
BUF_X1 \mifu/_458_ ( .A(\mifu/_015_ ), .Z(\mifu/_201_ ) );
BUF_X1 \mifu/_459_ ( .A(\mifu/_016_ ), .Z(\mifu/_202_ ) );
BUF_X1 \mifu/_460_ ( .A(\mifu/_017_ ), .Z(\mifu/_203_ ) );
BUF_X1 \mifu/_461_ ( .A(\mifu/_018_ ), .Z(\mifu/_204_ ) );
BUF_X1 \mifu/_462_ ( .A(\mifu/_019_ ), .Z(\mifu/_205_ ) );
BUF_X1 \mifu/_463_ ( .A(\mifu/_020_ ), .Z(\mifu/_206_ ) );
BUF_X1 \mifu/_464_ ( .A(\mifu/_021_ ), .Z(\mifu/_207_ ) );
BUF_X1 \mifu/_465_ ( .A(\mifu/_022_ ), .Z(\mifu/_208_ ) );
BUF_X1 \mifu/_466_ ( .A(\mifu/_023_ ), .Z(\mifu/_209_ ) );
BUF_X1 \mifu/_467_ ( .A(\mifu/_024_ ), .Z(\mifu/_210_ ) );
BUF_X1 \mifu/_468_ ( .A(\mifu/_025_ ), .Z(\mifu/_211_ ) );
BUF_X1 \mifu/_469_ ( .A(\mifu/_026_ ), .Z(\mifu/_212_ ) );
BUF_X1 \mifu/_470_ ( .A(\mifu/_027_ ), .Z(\mifu/_213_ ) );
BUF_X1 \mifu/_471_ ( .A(\mifu/_028_ ), .Z(\mifu/_214_ ) );
BUF_X1 \mifu/_472_ ( .A(\mifu/_029_ ), .Z(\mifu/_215_ ) );
BUF_X1 \mifu/_473_ ( .A(\mifu/_030_ ), .Z(\mifu/_216_ ) );
BUF_X1 \mifu/_474_ ( .A(\mifu/_031_ ), .Z(\mifu/_217_ ) );
BUF_X1 \mifu/_475_ ( .A(\mifu/_032_ ), .Z(\mifu/_218_ ) );
BUF_X1 \mifu/_476_ ( .A(\mifu/_033_ ), .Z(\mifu/_219_ ) );
BUF_X1 \mifu/_477_ ( .A(\mifu/_034_ ), .Z(\mifu/_220_ ) );
BUF_X1 \mifu/_478_ ( .A(\mifu/_035_ ), .Z(\mifu/_221_ ) );
BUF_X1 \mifu/_479_ ( .A(\mifu/_036_ ), .Z(\mifu/_222_ ) );
BUF_X1 \mifu/_480_ ( .A(\mifu/_037_ ), .Z(\mifu/_223_ ) );
INV_X32 \mlsu/_270_ ( .A(\mlsu/_193_ ), .ZN(\mlsu/_108_ ) );
NAND2_X1 \mlsu/_271_ ( .A1(\mlsu/_108_ ), .A2(\mlsu/_063_ ), .ZN(\mlsu/_109_ ) );
OR2_X1 \mlsu/_272_ ( .A1(\mlsu/_109_ ), .A2(\mlsu/_191_ ), .ZN(\mlsu/_110_ ) );
AOI22_X1 \mlsu/_273_ ( .A1(\mlsu/_191_ ), .A2(\mlsu/_105_ ), .B1(\mlsu/_193_ ), .B2(\mlsu/_106_ ), .ZN(\mlsu/_111_ ) );
AOI21_X1 \mlsu/_274_ ( .A(\mlsu/_072_ ), .B1(\mlsu/_110_ ), .B2(\mlsu/_111_ ), .ZN(\mlsu/_001_ ) );
NOR3_X4 \mlsu/_275_ ( .A1(\mlsu/_065_ ), .A2(\mlsu/_064_ ), .A3(\mlsu/_066_ ), .ZN(\mlsu/_112_ ) );
NAND2_X4 \mlsu/_276_ ( .A1(\mlsu/_112_ ), .A2(\mlsu/_188_ ), .ZN(\mlsu/_113_ ) );
BUF_X4 \mlsu/_277_ ( .A(\mlsu/_113_ ), .Z(\mlsu/_114_ ) );
OAI21_X1 \mlsu/_278_ ( .A(\mlsu/_024_ ), .B1(\mlsu/_065_ ), .B2(\mlsu/_064_ ), .ZN(\mlsu/_115_ ) );
NAND2_X1 \mlsu/_279_ ( .A1(\mlsu/_114_ ), .A2(\mlsu/_115_ ), .ZN(\mlsu/_189_ ) );
OAI21_X1 \mlsu/_280_ ( .A(\mlsu/_025_ ), .B1(\mlsu/_065_ ), .B2(\mlsu/_064_ ), .ZN(\mlsu/_116_ ) );
NAND2_X1 \mlsu/_281_ ( .A1(\mlsu/_114_ ), .A2(\mlsu/_116_ ), .ZN(\mlsu/_190_ ) );
OAI21_X1 \mlsu/_282_ ( .A(\mlsu/_002_ ), .B1(\mlsu/_065_ ), .B2(\mlsu/_064_ ), .ZN(\mlsu/_117_ ) );
NAND2_X1 \mlsu/_283_ ( .A1(\mlsu/_114_ ), .A2(\mlsu/_117_ ), .ZN(\mlsu/_160_ ) );
OAI21_X1 \mlsu/_284_ ( .A(\mlsu/_003_ ), .B1(\mlsu/_065_ ), .B2(\mlsu/_064_ ), .ZN(\mlsu/_118_ ) );
NAND2_X1 \mlsu/_285_ ( .A1(\mlsu/_114_ ), .A2(\mlsu/_118_ ), .ZN(\mlsu/_161_ ) );
OAI21_X1 \mlsu/_286_ ( .A(\mlsu/_004_ ), .B1(\mlsu/_065_ ), .B2(\mlsu/_064_ ), .ZN(\mlsu/_119_ ) );
NAND2_X1 \mlsu/_287_ ( .A1(\mlsu/_114_ ), .A2(\mlsu/_119_ ), .ZN(\mlsu/_162_ ) );
OAI21_X1 \mlsu/_288_ ( .A(\mlsu/_005_ ), .B1(\mlsu/_065_ ), .B2(\mlsu/_064_ ), .ZN(\mlsu/_120_ ) );
NAND2_X1 \mlsu/_289_ ( .A1(\mlsu/_114_ ), .A2(\mlsu/_120_ ), .ZN(\mlsu/_163_ ) );
OAI21_X1 \mlsu/_290_ ( .A(\mlsu/_006_ ), .B1(\mlsu/_065_ ), .B2(\mlsu/_064_ ), .ZN(\mlsu/_121_ ) );
NAND2_X1 \mlsu/_291_ ( .A1(\mlsu/_114_ ), .A2(\mlsu/_121_ ), .ZN(\mlsu/_164_ ) );
INV_X16 \mlsu/_292_ ( .A(\mlsu/_065_ ), .ZN(\mlsu/_122_ ) );
NAND2_X2 \mlsu/_293_ ( .A1(\mlsu/_122_ ), .A2(\mlsu/_064_ ), .ZN(\mlsu/_123_ ) );
INV_X2 \mlsu/_294_ ( .A(\mlsu/_007_ ), .ZN(\mlsu/_124_ ) );
OR3_X4 \mlsu/_295_ ( .A1(\mlsu/_123_ ), .A2(\mlsu/_066_ ), .A3(\mlsu/_124_ ), .ZN(\mlsu/_125_ ) );
AND2_X4 \mlsu/_296_ ( .A1(\mlsu/_125_ ), .A2(\mlsu/_113_ ), .ZN(\mlsu/_126_ ) );
NAND4_X1 \mlsu/_297_ ( .A1(\mlsu/_122_ ), .A2(\mlsu/_064_ ), .A3(\mlsu/_066_ ), .A4(\mlsu/_007_ ), .ZN(\mlsu/_127_ ) );
OAI211_X2 \mlsu/_298_ ( .A(\mlsu/_126_ ), .B(\mlsu/_127_ ), .C1(\mlsu/_122_ ), .C2(\mlsu/_124_ ), .ZN(\mlsu/_165_ ) );
BUF_X8 \mlsu/_299_ ( .A(\mlsu/_125_ ), .Z(\mlsu/_128_ ) );
NAND2_X1 \mlsu/_300_ ( .A1(\mlsu/_065_ ), .A2(\mlsu/_008_ ), .ZN(\mlsu/_129_ ) );
NAND3_X1 \mlsu/_301_ ( .A1(\mlsu/_128_ ), .A2(\mlsu/_114_ ), .A3(\mlsu/_129_ ), .ZN(\mlsu/_166_ ) );
NAND2_X1 \mlsu/_302_ ( .A1(\mlsu/_065_ ), .A2(\mlsu/_009_ ), .ZN(\mlsu/_130_ ) );
NAND3_X1 \mlsu/_303_ ( .A1(\mlsu/_128_ ), .A2(\mlsu/_114_ ), .A3(\mlsu/_130_ ), .ZN(\mlsu/_167_ ) );
NAND2_X1 \mlsu/_304_ ( .A1(\mlsu/_065_ ), .A2(\mlsu/_010_ ), .ZN(\mlsu/_131_ ) );
NAND3_X1 \mlsu/_305_ ( .A1(\mlsu/_128_ ), .A2(\mlsu/_114_ ), .A3(\mlsu/_131_ ), .ZN(\mlsu/_168_ ) );
BUF_X4 \mlsu/_306_ ( .A(\mlsu/_113_ ), .Z(\mlsu/_132_ ) );
NAND2_X1 \mlsu/_307_ ( .A1(\mlsu/_065_ ), .A2(\mlsu/_011_ ), .ZN(\mlsu/_133_ ) );
NAND3_X1 \mlsu/_308_ ( .A1(\mlsu/_128_ ), .A2(\mlsu/_132_ ), .A3(\mlsu/_133_ ), .ZN(\mlsu/_169_ ) );
NAND2_X1 \mlsu/_309_ ( .A1(\mlsu/_065_ ), .A2(\mlsu/_012_ ), .ZN(\mlsu/_134_ ) );
NAND3_X1 \mlsu/_310_ ( .A1(\mlsu/_128_ ), .A2(\mlsu/_132_ ), .A3(\mlsu/_134_ ), .ZN(\mlsu/_171_ ) );
NAND2_X1 \mlsu/_311_ ( .A1(\mlsu/_065_ ), .A2(\mlsu/_013_ ), .ZN(\mlsu/_135_ ) );
NAND3_X1 \mlsu/_312_ ( .A1(\mlsu/_128_ ), .A2(\mlsu/_132_ ), .A3(\mlsu/_135_ ), .ZN(\mlsu/_172_ ) );
NAND2_X1 \mlsu/_313_ ( .A1(\mlsu/_065_ ), .A2(\mlsu/_014_ ), .ZN(\mlsu/_136_ ) );
NAND3_X1 \mlsu/_314_ ( .A1(\mlsu/_128_ ), .A2(\mlsu/_132_ ), .A3(\mlsu/_136_ ), .ZN(\mlsu/_173_ ) );
NAND2_X1 \mlsu/_315_ ( .A1(\mlsu/_065_ ), .A2(\mlsu/_015_ ), .ZN(\mlsu/_137_ ) );
NAND3_X1 \mlsu/_316_ ( .A1(\mlsu/_128_ ), .A2(\mlsu/_132_ ), .A3(\mlsu/_137_ ), .ZN(\mlsu/_174_ ) );
NAND2_X1 \mlsu/_317_ ( .A1(\mlsu/_065_ ), .A2(\mlsu/_016_ ), .ZN(\mlsu/_138_ ) );
NAND3_X1 \mlsu/_318_ ( .A1(\mlsu/_128_ ), .A2(\mlsu/_132_ ), .A3(\mlsu/_138_ ), .ZN(\mlsu/_175_ ) );
NAND2_X1 \mlsu/_319_ ( .A1(\mlsu/_065_ ), .A2(\mlsu/_017_ ), .ZN(\mlsu/_139_ ) );
NAND3_X1 \mlsu/_320_ ( .A1(\mlsu/_128_ ), .A2(\mlsu/_132_ ), .A3(\mlsu/_139_ ), .ZN(\mlsu/_176_ ) );
NAND2_X1 \mlsu/_321_ ( .A1(\mlsu/_065_ ), .A2(\mlsu/_018_ ), .ZN(\mlsu/_140_ ) );
NAND3_X1 \mlsu/_322_ ( .A1(\mlsu/_125_ ), .A2(\mlsu/_132_ ), .A3(\mlsu/_140_ ), .ZN(\mlsu/_177_ ) );
NAND2_X1 \mlsu/_323_ ( .A1(\mlsu/_065_ ), .A2(\mlsu/_019_ ), .ZN(\mlsu/_141_ ) );
NAND3_X1 \mlsu/_324_ ( .A1(\mlsu/_125_ ), .A2(\mlsu/_132_ ), .A3(\mlsu/_141_ ), .ZN(\mlsu/_178_ ) );
NAND2_X1 \mlsu/_325_ ( .A1(\mlsu/_065_ ), .A2(\mlsu/_020_ ), .ZN(\mlsu/_142_ ) );
NAND3_X1 \mlsu/_326_ ( .A1(\mlsu/_125_ ), .A2(\mlsu/_132_ ), .A3(\mlsu/_142_ ), .ZN(\mlsu/_179_ ) );
NAND2_X1 \mlsu/_327_ ( .A1(\mlsu/_065_ ), .A2(\mlsu/_021_ ), .ZN(\mlsu/_143_ ) );
NAND3_X1 \mlsu/_328_ ( .A1(\mlsu/_125_ ), .A2(\mlsu/_113_ ), .A3(\mlsu/_143_ ), .ZN(\mlsu/_180_ ) );
NAND2_X1 \mlsu/_329_ ( .A1(\mlsu/_065_ ), .A2(\mlsu/_022_ ), .ZN(\mlsu/_144_ ) );
NAND3_X1 \mlsu/_330_ ( .A1(\mlsu/_125_ ), .A2(\mlsu/_113_ ), .A3(\mlsu/_144_ ), .ZN(\mlsu/_182_ ) );
NAND2_X1 \mlsu/_331_ ( .A1(\mlsu/_065_ ), .A2(\mlsu/_023_ ), .ZN(\mlsu/_145_ ) );
NAND3_X1 \mlsu/_332_ ( .A1(\mlsu/_125_ ), .A2(\mlsu/_113_ ), .A3(\mlsu/_145_ ), .ZN(\mlsu/_183_ ) );
NOR2_X4 \mlsu/_333_ ( .A1(\mlsu/_108_ ), .A2(\mlsu/_194_ ), .ZN(\mlsu/_146_ ) );
AND2_X4 \mlsu/_334_ ( .A1(\mlsu/_146_ ), .A2(\mlsu/_063_ ), .ZN(\mlsu/_147_ ) );
INV_X2 \mlsu/_335_ ( .A(\mlsu/_106_ ), .ZN(\mlsu/_148_ ) );
NOR2_X1 \mlsu/_336_ ( .A1(\mlsu/_146_ ), .A2(\mlsu/_148_ ), .ZN(\mlsu/_149_ ) );
NOR2_X2 \mlsu/_337_ ( .A1(\mlsu/_147_ ), .A2(\mlsu/_149_ ), .ZN(\mlsu/_150_ ) );
NOR2_X2 \mlsu/_338_ ( .A1(\mlsu/_150_ ), .A2(\mlsu/_192_ ), .ZN(\mlsu/_151_ ) );
MUX2_X1 \mlsu/_339_ ( .A(\mlsu/_107_ ), .B(\mlsu/_146_ ), .S(\mlsu/_151_ ), .Z(\mlsu/_030_ ) );
MUX2_X1 \mlsu/_340_ ( .A(\mlsu/_159_ ), .B(\mlsu/_073_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_031_ ) );
MUX2_X1 \mlsu/_341_ ( .A(\mlsu/_170_ ), .B(\mlsu/_084_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_032_ ) );
MUX2_X1 \mlsu/_342_ ( .A(\mlsu/_181_ ), .B(\mlsu/_095_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_033_ ) );
MUX2_X1 \mlsu/_343_ ( .A(\mlsu/_184_ ), .B(\mlsu/_098_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_034_ ) );
MUX2_X1 \mlsu/_344_ ( .A(\mlsu/_185_ ), .B(\mlsu/_099_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_035_ ) );
MUX2_X1 \mlsu/_345_ ( .A(\mlsu/_186_ ), .B(\mlsu/_100_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_036_ ) );
MUX2_X1 \mlsu/_346_ ( .A(\mlsu/_187_ ), .B(\mlsu/_101_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_037_ ) );
MUX2_X1 \mlsu/_347_ ( .A(\mlsu/_188_ ), .B(\mlsu/_102_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_038_ ) );
MUX2_X1 \mlsu/_348_ ( .A(\mlsu/_024_ ), .B(\mlsu/_103_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_039_ ) );
MUX2_X1 \mlsu/_349_ ( .A(\mlsu/_025_ ), .B(\mlsu/_104_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_040_ ) );
MUX2_X1 \mlsu/_350_ ( .A(\mlsu/_002_ ), .B(\mlsu/_074_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_041_ ) );
MUX2_X1 \mlsu/_351_ ( .A(\mlsu/_003_ ), .B(\mlsu/_075_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_042_ ) );
MUX2_X1 \mlsu/_352_ ( .A(\mlsu/_004_ ), .B(\mlsu/_076_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_043_ ) );
MUX2_X1 \mlsu/_353_ ( .A(\mlsu/_005_ ), .B(\mlsu/_077_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_044_ ) );
MUX2_X1 \mlsu/_354_ ( .A(\mlsu/_006_ ), .B(\mlsu/_078_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_045_ ) );
MUX2_X1 \mlsu/_355_ ( .A(\mlsu/_007_ ), .B(\mlsu/_079_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_046_ ) );
MUX2_X1 \mlsu/_356_ ( .A(\mlsu/_008_ ), .B(\mlsu/_080_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_047_ ) );
MUX2_X1 \mlsu/_357_ ( .A(\mlsu/_009_ ), .B(\mlsu/_081_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_048_ ) );
MUX2_X1 \mlsu/_358_ ( .A(\mlsu/_010_ ), .B(\mlsu/_082_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_049_ ) );
MUX2_X1 \mlsu/_359_ ( .A(\mlsu/_011_ ), .B(\mlsu/_083_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_050_ ) );
MUX2_X1 \mlsu/_360_ ( .A(\mlsu/_012_ ), .B(\mlsu/_085_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_051_ ) );
MUX2_X1 \mlsu/_361_ ( .A(\mlsu/_013_ ), .B(\mlsu/_086_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_052_ ) );
MUX2_X1 \mlsu/_362_ ( .A(\mlsu/_014_ ), .B(\mlsu/_087_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_053_ ) );
MUX2_X1 \mlsu/_363_ ( .A(\mlsu/_015_ ), .B(\mlsu/_088_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_054_ ) );
MUX2_X1 \mlsu/_364_ ( .A(\mlsu/_016_ ), .B(\mlsu/_089_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_055_ ) );
MUX2_X1 \mlsu/_365_ ( .A(\mlsu/_017_ ), .B(\mlsu/_090_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_056_ ) );
MUX2_X1 \mlsu/_366_ ( .A(\mlsu/_018_ ), .B(\mlsu/_091_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_057_ ) );
MUX2_X1 \mlsu/_367_ ( .A(\mlsu/_019_ ), .B(\mlsu/_092_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_058_ ) );
MUX2_X1 \mlsu/_368_ ( .A(\mlsu/_020_ ), .B(\mlsu/_093_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_059_ ) );
MUX2_X1 \mlsu/_369_ ( .A(\mlsu/_021_ ), .B(\mlsu/_094_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_060_ ) );
MUX2_X1 \mlsu/_370_ ( .A(\mlsu/_022_ ), .B(\mlsu/_096_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_061_ ) );
MUX2_X1 \mlsu/_371_ ( .A(\mlsu/_023_ ), .B(\mlsu/_097_ ), .S(\mlsu/_105_ ), .Z(\mlsu/_062_ ) );
OR3_X4 \mlsu/_372_ ( .A1(\mlsu/_108_ ), .A2(\mlsu/_194_ ), .A3(\mlsu/_063_ ), .ZN(\mlsu/_152_ ) );
NAND3_X2 \mlsu/_373_ ( .A1(\mlsu/_152_ ), .A2(\mlsu/_069_ ), .A3(\mlsu/_070_ ), .ZN(\mlsu/_153_ ) );
NAND3_X1 \mlsu/_374_ ( .A1(\mlsu/_150_ ), .A2(\mlsu/_153_ ), .A3(\mlsu/_070_ ), .ZN(\mlsu/_154_ ) );
INV_X1 \mlsu/_375_ ( .A(\mlsu/_147_ ), .ZN(\mlsu/_155_ ) );
AOI21_X1 \mlsu/_376_ ( .A(\mlsu/_192_ ), .B1(\mlsu/_154_ ), .B2(\mlsu/_155_ ), .ZN(\mlsu/_026_ ) );
NAND4_X1 \mlsu/_377_ ( .A1(\mlsu/_148_ ), .A2(\mlsu/_069_ ), .A3(\mlsu/_070_ ), .A4(\mlsu/_071_ ), .ZN(\mlsu/_156_ ) );
AOI211_X2 \mlsu/_378_ ( .A(\mlsu/_192_ ), .B(\mlsu/_146_ ), .C1(\mlsu/_148_ ), .C2(\mlsu/_156_ ), .ZN(\mlsu/_027_ ) );
NAND2_X1 \mlsu/_379_ ( .A1(\mlsu/_148_ ), .A2(\mlsu/_194_ ), .ZN(\mlsu/_157_ ) );
AOI21_X1 \mlsu/_380_ ( .A(\mlsu/_192_ ), .B1(\mlsu/_155_ ), .B2(\mlsu/_157_ ), .ZN(\mlsu/_028_ ) );
AOI21_X1 \mlsu/_381_ ( .A(\mlsu/_068_ ), .B1(\mlsu/_191_ ), .B2(\mlsu/_063_ ), .ZN(\mlsu/_158_ ) );
AOI211_X2 \mlsu/_382_ ( .A(\mlsu/_192_ ), .B(\mlsu/_158_ ), .C1(\mlsu/_068_ ), .C2(\mlsu/_067_ ), .ZN(\mlsu/_029_ ) );
DFF_X1 \mlsu/_383_ ( .CK(clk ), .D(\mlsu/_000_ ), .Q(lsu_finish ), .QN(\mlsu/_232_ ) );
DFF_X1 \mlsu/_384_ ( .CK(clk ), .D(\mlsu/_233_ ), .Q(lsu_awvalid ), .QN(\mlsu/_231_ ) );
DFF_X1 \mlsu/_385_ ( .CK(clk ), .D(\mlsu/_234_ ), .Q(lsu_bready ), .QN(\mlsu/_230_ ) );
DFF_X1 \mlsu/_386_ ( .CK(clk ), .D(\mlsu/_235_ ), .Q(\mlsu/write_wait_ready ), .QN(\mlsu/_229_ ) );
DFF_X1 \mlsu/_387_ ( .CK(clk ), .D(\mlsu/_236_ ), .Q(lsu_arvalid ), .QN(\mlsu/_228_ ) );
DFF_X1 \mlsu/_388_ ( .CK(clk ), .D(\mlsu/_237_ ), .Q(lsu_wvalid ), .QN(\mlsu/_227_ ) );
DFF_X1 \mlsu/_389_ ( .CK(clk ), .D(\mlsu/_238_ ), .Q(\mem_rdata[0] ), .QN(\mlsu/_226_ ) );
DFF_X1 \mlsu/_390_ ( .CK(clk ), .D(\mlsu/_239_ ), .Q(\mem_rdata[1] ), .QN(\mlsu/_225_ ) );
DFF_X1 \mlsu/_391_ ( .CK(clk ), .D(\mlsu/_240_ ), .Q(\mem_rdata[2] ), .QN(\mlsu/_224_ ) );
DFF_X1 \mlsu/_392_ ( .CK(clk ), .D(\mlsu/_241_ ), .Q(\mem_rdata[3] ), .QN(\mlsu/_223_ ) );
DFF_X1 \mlsu/_393_ ( .CK(clk ), .D(\mlsu/_242_ ), .Q(\mem_rdata[4] ), .QN(\mlsu/_222_ ) );
DFF_X1 \mlsu/_394_ ( .CK(clk ), .D(\mlsu/_243_ ), .Q(\mem_rdata[5] ), .QN(\mlsu/_221_ ) );
DFF_X1 \mlsu/_395_ ( .CK(clk ), .D(\mlsu/_244_ ), .Q(\mem_rdata[6] ), .QN(\mlsu/_220_ ) );
DFF_X1 \mlsu/_396_ ( .CK(clk ), .D(\mlsu/_245_ ), .Q(\mem_rdata[7] ), .QN(\mlsu/_219_ ) );
DFF_X1 \mlsu/_397_ ( .CK(clk ), .D(\mlsu/_246_ ), .Q(\mlsu/_rdata[8] ), .QN(\mlsu/_218_ ) );
DFF_X1 \mlsu/_398_ ( .CK(clk ), .D(\mlsu/_247_ ), .Q(\mlsu/_rdata[9] ), .QN(\mlsu/_217_ ) );
DFF_X1 \mlsu/_399_ ( .CK(clk ), .D(\mlsu/_248_ ), .Q(\mlsu/_rdata[10] ), .QN(\mlsu/_216_ ) );
DFF_X1 \mlsu/_400_ ( .CK(clk ), .D(\mlsu/_249_ ), .Q(\mlsu/_rdata[11] ), .QN(\mlsu/_215_ ) );
DFF_X1 \mlsu/_401_ ( .CK(clk ), .D(\mlsu/_250_ ), .Q(\mlsu/_rdata[12] ), .QN(\mlsu/_214_ ) );
DFF_X1 \mlsu/_402_ ( .CK(clk ), .D(\mlsu/_251_ ), .Q(\mlsu/_rdata[13] ), .QN(\mlsu/_213_ ) );
DFF_X1 \mlsu/_403_ ( .CK(clk ), .D(\mlsu/_252_ ), .Q(\mlsu/_rdata[14] ), .QN(\mlsu/_212_ ) );
DFF_X1 \mlsu/_404_ ( .CK(clk ), .D(\mlsu/_253_ ), .Q(\mlsu/_rdata[15] ), .QN(\mlsu/_211_ ) );
DFF_X1 \mlsu/_405_ ( .CK(clk ), .D(\mlsu/_254_ ), .Q(\mlsu/_rdata[16] ), .QN(\mlsu/_210_ ) );
DFF_X1 \mlsu/_406_ ( .CK(clk ), .D(\mlsu/_255_ ), .Q(\mlsu/_rdata[17] ), .QN(\mlsu/_209_ ) );
DFF_X1 \mlsu/_407_ ( .CK(clk ), .D(\mlsu/_256_ ), .Q(\mlsu/_rdata[18] ), .QN(\mlsu/_208_ ) );
DFF_X1 \mlsu/_408_ ( .CK(clk ), .D(\mlsu/_257_ ), .Q(\mlsu/_rdata[19] ), .QN(\mlsu/_207_ ) );
DFF_X1 \mlsu/_409_ ( .CK(clk ), .D(\mlsu/_258_ ), .Q(\mlsu/_rdata[20] ), .QN(\mlsu/_206_ ) );
DFF_X1 \mlsu/_410_ ( .CK(clk ), .D(\mlsu/_259_ ), .Q(\mlsu/_rdata[21] ), .QN(\mlsu/_205_ ) );
DFF_X1 \mlsu/_411_ ( .CK(clk ), .D(\mlsu/_260_ ), .Q(\mlsu/_rdata[22] ), .QN(\mlsu/_204_ ) );
DFF_X1 \mlsu/_412_ ( .CK(clk ), .D(\mlsu/_261_ ), .Q(\mlsu/_rdata[23] ), .QN(\mlsu/_203_ ) );
DFF_X1 \mlsu/_413_ ( .CK(clk ), .D(\mlsu/_262_ ), .Q(\mlsu/_rdata[24] ), .QN(\mlsu/_202_ ) );
DFF_X1 \mlsu/_414_ ( .CK(clk ), .D(\mlsu/_263_ ), .Q(\mlsu/_rdata[25] ), .QN(\mlsu/_201_ ) );
DFF_X1 \mlsu/_415_ ( .CK(clk ), .D(\mlsu/_264_ ), .Q(\mlsu/_rdata[26] ), .QN(\mlsu/_200_ ) );
DFF_X1 \mlsu/_416_ ( .CK(clk ), .D(\mlsu/_265_ ), .Q(\mlsu/_rdata[27] ), .QN(\mlsu/_199_ ) );
DFF_X1 \mlsu/_417_ ( .CK(clk ), .D(\mlsu/_266_ ), .Q(\mlsu/_rdata[28] ), .QN(\mlsu/_198_ ) );
DFF_X1 \mlsu/_418_ ( .CK(clk ), .D(\mlsu/_267_ ), .Q(\mlsu/_rdata[29] ), .QN(\mlsu/_197_ ) );
DFF_X1 \mlsu/_419_ ( .CK(clk ), .D(\mlsu/_268_ ), .Q(\mlsu/_rdata[30] ), .QN(\mlsu/_196_ ) );
DFF_X1 \mlsu/_420_ ( .CK(clk ), .D(\mlsu/_269_ ), .Q(\mlsu/_rdata[31] ), .QN(\mlsu/_195_ ) );
BUF_X1 \mlsu/_421_ ( .A(\mem_rdata[0] ), .Z(\mlsu/_rdata[0] ) );
BUF_X1 \mlsu/_422_ ( .A(\mem_rdata[1] ), .Z(\mlsu/_rdata[1] ) );
BUF_X1 \mlsu/_423_ ( .A(\mem_rdata[2] ), .Z(\mlsu/_rdata[2] ) );
BUF_X1 \mlsu/_424_ ( .A(\mem_rdata[3] ), .Z(\mlsu/_rdata[3] ) );
BUF_X1 \mlsu/_425_ ( .A(\mem_rdata[4] ), .Z(\mlsu/_rdata[4] ) );
BUF_X1 \mlsu/_426_ ( .A(\mem_rdata[5] ), .Z(\mlsu/_rdata[5] ) );
BUF_X1 \mlsu/_427_ ( .A(\mem_rdata[6] ), .Z(\mlsu/_rdata[6] ) );
BUF_X1 \mlsu/_428_ ( .A(\mem_rdata[7] ), .Z(\mlsu/_rdata[7] ) );
BUF_X1 \mlsu/_429_ ( .A(\alu_result[0] ), .Z(\lsu_araddr[0] ) );
BUF_X1 \mlsu/_430_ ( .A(\alu_result[1] ), .Z(\lsu_araddr[1] ) );
BUF_X1 \mlsu/_431_ ( .A(\alu_result[2] ), .Z(\lsu_araddr[2] ) );
BUF_X1 \mlsu/_432_ ( .A(\alu_result[3] ), .Z(\lsu_araddr[3] ) );
BUF_X1 \mlsu/_433_ ( .A(\alu_result[4] ), .Z(\lsu_araddr[4] ) );
BUF_X1 \mlsu/_434_ ( .A(\alu_result[5] ), .Z(\lsu_araddr[5] ) );
BUF_X1 \mlsu/_435_ ( .A(\alu_result[6] ), .Z(\lsu_araddr[6] ) );
BUF_X1 \mlsu/_436_ ( .A(\alu_result[7] ), .Z(\lsu_araddr[7] ) );
BUF_X1 \mlsu/_437_ ( .A(\alu_result[8] ), .Z(\lsu_araddr[8] ) );
BUF_X1 \mlsu/_438_ ( .A(\alu_result[9] ), .Z(\lsu_araddr[9] ) );
BUF_X1 \mlsu/_439_ ( .A(\alu_result[10] ), .Z(\lsu_araddr[10] ) );
BUF_X1 \mlsu/_440_ ( .A(\alu_result[11] ), .Z(\lsu_araddr[11] ) );
BUF_X1 \mlsu/_441_ ( .A(\alu_result[12] ), .Z(\lsu_araddr[12] ) );
BUF_X1 \mlsu/_442_ ( .A(\alu_result[13] ), .Z(\lsu_araddr[13] ) );
BUF_X1 \mlsu/_443_ ( .A(\alu_result[14] ), .Z(\lsu_araddr[14] ) );
BUF_X1 \mlsu/_444_ ( .A(\alu_result[15] ), .Z(\lsu_araddr[15] ) );
BUF_X1 \mlsu/_445_ ( .A(\alu_result[16] ), .Z(\lsu_araddr[16] ) );
BUF_X1 \mlsu/_446_ ( .A(\alu_result[17] ), .Z(\lsu_araddr[17] ) );
BUF_X1 \mlsu/_447_ ( .A(\alu_result[18] ), .Z(\lsu_araddr[18] ) );
BUF_X1 \mlsu/_448_ ( .A(\alu_result[19] ), .Z(\lsu_araddr[19] ) );
BUF_X1 \mlsu/_449_ ( .A(\alu_result[20] ), .Z(\lsu_araddr[20] ) );
BUF_X1 \mlsu/_450_ ( .A(\alu_result[21] ), .Z(\lsu_araddr[21] ) );
BUF_X1 \mlsu/_451_ ( .A(\alu_result[22] ), .Z(\lsu_araddr[22] ) );
BUF_X1 \mlsu/_452_ ( .A(\alu_result[23] ), .Z(\lsu_araddr[23] ) );
BUF_X1 \mlsu/_453_ ( .A(\alu_result[24] ), .Z(\lsu_araddr[24] ) );
BUF_X1 \mlsu/_454_ ( .A(\alu_result[25] ), .Z(\lsu_araddr[25] ) );
BUF_X1 \mlsu/_455_ ( .A(\alu_result[26] ), .Z(\lsu_araddr[26] ) );
BUF_X1 \mlsu/_456_ ( .A(\alu_result[27] ), .Z(\lsu_araddr[27] ) );
BUF_X1 \mlsu/_457_ ( .A(\alu_result[28] ), .Z(\lsu_araddr[28] ) );
BUF_X1 \mlsu/_458_ ( .A(\alu_result[29] ), .Z(\lsu_araddr[29] ) );
BUF_X1 \mlsu/_459_ ( .A(\alu_result[30] ), .Z(\lsu_araddr[30] ) );
BUF_X1 \mlsu/_460_ ( .A(\alu_result[31] ), .Z(\lsu_araddr[31] ) );
BUF_X1 \mlsu/_461_ ( .A(\alu_result[0] ), .Z(\lsu_awaddr[0] ) );
BUF_X1 \mlsu/_462_ ( .A(\alu_result[1] ), .Z(\lsu_awaddr[1] ) );
BUF_X1 \mlsu/_463_ ( .A(\alu_result[2] ), .Z(\lsu_awaddr[2] ) );
BUF_X1 \mlsu/_464_ ( .A(\alu_result[3] ), .Z(\lsu_awaddr[3] ) );
BUF_X1 \mlsu/_465_ ( .A(\alu_result[4] ), .Z(\lsu_awaddr[4] ) );
BUF_X1 \mlsu/_466_ ( .A(\alu_result[5] ), .Z(\lsu_awaddr[5] ) );
BUF_X1 \mlsu/_467_ ( .A(\alu_result[6] ), .Z(\lsu_awaddr[6] ) );
BUF_X1 \mlsu/_468_ ( .A(\alu_result[7] ), .Z(\lsu_awaddr[7] ) );
BUF_X1 \mlsu/_469_ ( .A(\alu_result[8] ), .Z(\lsu_awaddr[8] ) );
BUF_X1 \mlsu/_470_ ( .A(\alu_result[9] ), .Z(\lsu_awaddr[9] ) );
BUF_X1 \mlsu/_471_ ( .A(\alu_result[10] ), .Z(\lsu_awaddr[10] ) );
BUF_X1 \mlsu/_472_ ( .A(\alu_result[11] ), .Z(\lsu_awaddr[11] ) );
BUF_X1 \mlsu/_473_ ( .A(\alu_result[12] ), .Z(\lsu_awaddr[12] ) );
BUF_X1 \mlsu/_474_ ( .A(\alu_result[13] ), .Z(\lsu_awaddr[13] ) );
BUF_X1 \mlsu/_475_ ( .A(\alu_result[14] ), .Z(\lsu_awaddr[14] ) );
BUF_X1 \mlsu/_476_ ( .A(\alu_result[15] ), .Z(\lsu_awaddr[15] ) );
BUF_X1 \mlsu/_477_ ( .A(\alu_result[16] ), .Z(\lsu_awaddr[16] ) );
BUF_X1 \mlsu/_478_ ( .A(\alu_result[17] ), .Z(\lsu_awaddr[17] ) );
BUF_X1 \mlsu/_479_ ( .A(\alu_result[18] ), .Z(\lsu_awaddr[18] ) );
BUF_X1 \mlsu/_480_ ( .A(\alu_result[19] ), .Z(\lsu_awaddr[19] ) );
BUF_X1 \mlsu/_481_ ( .A(\alu_result[20] ), .Z(\lsu_awaddr[20] ) );
BUF_X1 \mlsu/_482_ ( .A(\alu_result[21] ), .Z(\lsu_awaddr[21] ) );
BUF_X1 \mlsu/_483_ ( .A(\alu_result[22] ), .Z(\lsu_awaddr[22] ) );
BUF_X1 \mlsu/_484_ ( .A(\alu_result[23] ), .Z(\lsu_awaddr[23] ) );
BUF_X1 \mlsu/_485_ ( .A(\alu_result[24] ), .Z(\lsu_awaddr[24] ) );
BUF_X1 \mlsu/_486_ ( .A(\alu_result[25] ), .Z(\lsu_awaddr[25] ) );
BUF_X1 \mlsu/_487_ ( .A(\alu_result[26] ), .Z(\lsu_awaddr[26] ) );
BUF_X1 \mlsu/_488_ ( .A(\alu_result[27] ), .Z(\lsu_awaddr[27] ) );
BUF_X1 \mlsu/_489_ ( .A(\alu_result[28] ), .Z(\lsu_awaddr[28] ) );
BUF_X1 \mlsu/_490_ ( .A(\alu_result[29] ), .Z(\lsu_awaddr[29] ) );
BUF_X1 \mlsu/_491_ ( .A(\alu_result[30] ), .Z(\lsu_awaddr[30] ) );
BUF_X1 \mlsu/_492_ ( .A(\alu_result[31] ), .Z(\lsu_awaddr[31] ) );
BUF_X1 \mlsu/_493_ ( .A(1'b0 ), .Z(lsu_rready ) );
BUF_X1 \mlsu/_494_ ( .A(\mem_wdata[0] ), .Z(\lsu_wdata[0] ) );
BUF_X1 \mlsu/_495_ ( .A(\mem_wdata[1] ), .Z(\lsu_wdata[1] ) );
BUF_X1 \mlsu/_496_ ( .A(\mem_wdata[2] ), .Z(\lsu_wdata[2] ) );
BUF_X1 \mlsu/_497_ ( .A(\mem_wdata[3] ), .Z(\lsu_wdata[3] ) );
BUF_X1 \mlsu/_498_ ( .A(\mem_wdata[4] ), .Z(\lsu_wdata[4] ) );
BUF_X1 \mlsu/_499_ ( .A(\mem_wdata[5] ), .Z(\lsu_wdata[5] ) );
BUF_X1 \mlsu/_500_ ( .A(\mem_wdata[6] ), .Z(\lsu_wdata[6] ) );
BUF_X1 \mlsu/_501_ ( .A(\mem_wdata[7] ), .Z(\lsu_wdata[7] ) );
BUF_X1 \mlsu/_502_ ( .A(\mem_wdata[8] ), .Z(\lsu_wdata[8] ) );
BUF_X1 \mlsu/_503_ ( .A(\mem_wdata[9] ), .Z(\lsu_wdata[9] ) );
BUF_X1 \mlsu/_504_ ( .A(\mem_wdata[10] ), .Z(\lsu_wdata[10] ) );
BUF_X1 \mlsu/_505_ ( .A(\mem_wdata[11] ), .Z(\lsu_wdata[11] ) );
BUF_X1 \mlsu/_506_ ( .A(\mem_wdata[12] ), .Z(\lsu_wdata[12] ) );
BUF_X1 \mlsu/_507_ ( .A(\mem_wdata[13] ), .Z(\lsu_wdata[13] ) );
BUF_X1 \mlsu/_508_ ( .A(\mem_wdata[14] ), .Z(\lsu_wdata[14] ) );
BUF_X1 \mlsu/_509_ ( .A(\mem_wdata[15] ), .Z(\lsu_wdata[15] ) );
BUF_X1 \mlsu/_510_ ( .A(\mem_wdata[16] ), .Z(\lsu_wdata[16] ) );
BUF_X1 \mlsu/_511_ ( .A(\mem_wdata[17] ), .Z(\lsu_wdata[17] ) );
BUF_X1 \mlsu/_512_ ( .A(\mem_wdata[18] ), .Z(\lsu_wdata[18] ) );
BUF_X1 \mlsu/_513_ ( .A(\mem_wdata[19] ), .Z(\lsu_wdata[19] ) );
BUF_X1 \mlsu/_514_ ( .A(\mem_wdata[20] ), .Z(\lsu_wdata[20] ) );
BUF_X1 \mlsu/_515_ ( .A(\mem_wdata[21] ), .Z(\lsu_wdata[21] ) );
BUF_X1 \mlsu/_516_ ( .A(\mem_wdata[22] ), .Z(\lsu_wdata[22] ) );
BUF_X1 \mlsu/_517_ ( .A(\mem_wdata[23] ), .Z(\lsu_wdata[23] ) );
BUF_X1 \mlsu/_518_ ( .A(\mem_wdata[24] ), .Z(\lsu_wdata[24] ) );
BUF_X1 \mlsu/_519_ ( .A(\mem_wdata[25] ), .Z(\lsu_wdata[25] ) );
BUF_X1 \mlsu/_520_ ( .A(\mem_wdata[26] ), .Z(\lsu_wdata[26] ) );
BUF_X1 \mlsu/_521_ ( .A(\mem_wdata[27] ), .Z(\lsu_wdata[27] ) );
BUF_X1 \mlsu/_522_ ( .A(\mem_wdata[28] ), .Z(\lsu_wdata[28] ) );
BUF_X1 \mlsu/_523_ ( .A(\mem_wdata[29] ), .Z(\lsu_wdata[29] ) );
BUF_X1 \mlsu/_524_ ( .A(\mem_wdata[30] ), .Z(\lsu_wdata[30] ) );
BUF_X1 \mlsu/_525_ ( .A(\mem_wdata[31] ), .Z(\lsu_wdata[31] ) );
BUF_X1 \mlsu/_526_ ( .A(\wmask[0] ), .Z(\lsu_wstrb[0] ) );
BUF_X1 \mlsu/_527_ ( .A(\wmask[1] ), .Z(\lsu_wstrb[1] ) );
BUF_X1 \mlsu/_528_ ( .A(\wmask[2] ), .Z(\lsu_wstrb[2] ) );
BUF_X1 \mlsu/_529_ ( .A(\wmask[3] ), .Z(\lsu_wstrb[3] ) );
BUF_X1 \mlsu/_530_ ( .A(\wmask[4] ), .Z(\lsu_wstrb[4] ) );
BUF_X1 \mlsu/_531_ ( .A(\wmask[5] ), .Z(\lsu_wstrb[5] ) );
BUF_X1 \mlsu/_532_ ( .A(\wmask[6] ), .Z(\lsu_wstrb[6] ) );
BUF_X1 \mlsu/_533_ ( .A(\wmask[7] ), .Z(\lsu_wstrb[7] ) );
BUF_X1 \mlsu/_534_ ( .A(mem_ren ), .Z(\mlsu/_191_ ) );
BUF_X1 \mlsu/_535_ ( .A(lsu_arvalid ), .Z(\mlsu/_068_ ) );
BUF_X1 \mlsu/_536_ ( .A(mem_wen ), .Z(\mlsu/_193_ ) );
BUF_X1 \mlsu/_537_ ( .A(\mlsu/write_wait_ready ), .Z(\mlsu/_194_ ) );
BUF_X1 \mlsu/_538_ ( .A(lsu_arready ), .Z(\mlsu/_067_ ) );
BUF_X1 \mlsu/_539_ ( .A(inst_valid ), .Z(\mlsu/_063_ ) );
BUF_X1 \mlsu/_540_ ( .A(rst ), .Z(\mlsu/_192_ ) );
BUF_X1 \mlsu/_541_ ( .A(lsu_awready ), .Z(\mlsu/_069_ ) );
BUF_X1 \mlsu/_542_ ( .A(lsu_awvalid ), .Z(\mlsu/_070_ ) );
BUF_X1 \mlsu/_543_ ( .A(lsu_wready ), .Z(\mlsu/_106_ ) );
BUF_X1 \mlsu/_544_ ( .A(lsu_rvalid ), .Z(\mlsu/_105_ ) );
BUF_X1 \mlsu/_545_ ( .A(lsu_finish ), .Z(\mlsu/_072_ ) );
BUF_X1 \mlsu/_546_ ( .A(\mlsu/_001_ ), .Z(\mlsu/_000_ ) );
BUF_X1 \mlsu/_547_ ( .A(\load_ctl[1] ), .Z(\mlsu/_065_ ) );
BUF_X1 \mlsu/_548_ ( .A(\load_ctl[0] ), .Z(\mlsu/_064_ ) );
BUF_X1 \mlsu/_549_ ( .A(\load_ctl[2] ), .Z(\mlsu/_066_ ) );
BUF_X1 \mlsu/_550_ ( .A(\mlsu/_rdata[8] ), .Z(\mlsu/_024_ ) );
BUF_X1 \mlsu/_551_ ( .A(\mem_rdata[7] ), .Z(\mlsu/_188_ ) );
BUF_X1 \mlsu/_552_ ( .A(\mlsu/_189_ ), .Z(\mem_rdata[8] ) );
BUF_X1 \mlsu/_553_ ( .A(\mlsu/_rdata[9] ), .Z(\mlsu/_025_ ) );
BUF_X1 \mlsu/_554_ ( .A(\mlsu/_190_ ), .Z(\mem_rdata[9] ) );
BUF_X1 \mlsu/_555_ ( .A(\mlsu/_rdata[10] ), .Z(\mlsu/_002_ ) );
BUF_X1 \mlsu/_556_ ( .A(\mlsu/_160_ ), .Z(\mem_rdata[10] ) );
BUF_X1 \mlsu/_557_ ( .A(\mlsu/_rdata[11] ), .Z(\mlsu/_003_ ) );
BUF_X1 \mlsu/_558_ ( .A(\mlsu/_161_ ), .Z(\mem_rdata[11] ) );
BUF_X1 \mlsu/_559_ ( .A(\mlsu/_rdata[12] ), .Z(\mlsu/_004_ ) );
BUF_X1 \mlsu/_560_ ( .A(\mlsu/_162_ ), .Z(\mem_rdata[12] ) );
BUF_X1 \mlsu/_561_ ( .A(\mlsu/_rdata[13] ), .Z(\mlsu/_005_ ) );
BUF_X1 \mlsu/_562_ ( .A(\mlsu/_163_ ), .Z(\mem_rdata[13] ) );
BUF_X1 \mlsu/_563_ ( .A(\mlsu/_rdata[14] ), .Z(\mlsu/_006_ ) );
BUF_X1 \mlsu/_564_ ( .A(\mlsu/_164_ ), .Z(\mem_rdata[14] ) );
BUF_X1 \mlsu/_565_ ( .A(\mlsu/_rdata[15] ), .Z(\mlsu/_007_ ) );
BUF_X1 \mlsu/_566_ ( .A(\mlsu/_165_ ), .Z(\mem_rdata[15] ) );
BUF_X1 \mlsu/_567_ ( .A(\mlsu/_rdata[16] ), .Z(\mlsu/_008_ ) );
BUF_X1 \mlsu/_568_ ( .A(\mlsu/_166_ ), .Z(\mem_rdata[16] ) );
BUF_X1 \mlsu/_569_ ( .A(\mlsu/_rdata[17] ), .Z(\mlsu/_009_ ) );
BUF_X1 \mlsu/_570_ ( .A(\mlsu/_167_ ), .Z(\mem_rdata[17] ) );
BUF_X1 \mlsu/_571_ ( .A(\mlsu/_rdata[18] ), .Z(\mlsu/_010_ ) );
BUF_X1 \mlsu/_572_ ( .A(\mlsu/_168_ ), .Z(\mem_rdata[18] ) );
BUF_X1 \mlsu/_573_ ( .A(\mlsu/_rdata[19] ), .Z(\mlsu/_011_ ) );
BUF_X1 \mlsu/_574_ ( .A(\mlsu/_169_ ), .Z(\mem_rdata[19] ) );
BUF_X1 \mlsu/_575_ ( .A(\mlsu/_rdata[20] ), .Z(\mlsu/_012_ ) );
BUF_X1 \mlsu/_576_ ( .A(\mlsu/_171_ ), .Z(\mem_rdata[20] ) );
BUF_X1 \mlsu/_577_ ( .A(\mlsu/_rdata[21] ), .Z(\mlsu/_013_ ) );
BUF_X1 \mlsu/_578_ ( .A(\mlsu/_172_ ), .Z(\mem_rdata[21] ) );
BUF_X1 \mlsu/_579_ ( .A(\mlsu/_rdata[22] ), .Z(\mlsu/_014_ ) );
BUF_X1 \mlsu/_580_ ( .A(\mlsu/_173_ ), .Z(\mem_rdata[22] ) );
BUF_X1 \mlsu/_581_ ( .A(\mlsu/_rdata[23] ), .Z(\mlsu/_015_ ) );
BUF_X1 \mlsu/_582_ ( .A(\mlsu/_174_ ), .Z(\mem_rdata[23] ) );
BUF_X1 \mlsu/_583_ ( .A(\mlsu/_rdata[24] ), .Z(\mlsu/_016_ ) );
BUF_X1 \mlsu/_584_ ( .A(\mlsu/_175_ ), .Z(\mem_rdata[24] ) );
BUF_X1 \mlsu/_585_ ( .A(\mlsu/_rdata[25] ), .Z(\mlsu/_017_ ) );
BUF_X1 \mlsu/_586_ ( .A(\mlsu/_176_ ), .Z(\mem_rdata[25] ) );
BUF_X1 \mlsu/_587_ ( .A(\mlsu/_rdata[26] ), .Z(\mlsu/_018_ ) );
BUF_X1 \mlsu/_588_ ( .A(\mlsu/_177_ ), .Z(\mem_rdata[26] ) );
BUF_X1 \mlsu/_589_ ( .A(\mlsu/_rdata[27] ), .Z(\mlsu/_019_ ) );
BUF_X1 \mlsu/_590_ ( .A(\mlsu/_178_ ), .Z(\mem_rdata[27] ) );
BUF_X1 \mlsu/_591_ ( .A(\mlsu/_rdata[28] ), .Z(\mlsu/_020_ ) );
BUF_X1 \mlsu/_592_ ( .A(\mlsu/_179_ ), .Z(\mem_rdata[28] ) );
BUF_X1 \mlsu/_593_ ( .A(\mlsu/_rdata[29] ), .Z(\mlsu/_021_ ) );
BUF_X1 \mlsu/_594_ ( .A(\mlsu/_180_ ), .Z(\mem_rdata[29] ) );
BUF_X1 \mlsu/_595_ ( .A(\mlsu/_rdata[30] ), .Z(\mlsu/_022_ ) );
BUF_X1 \mlsu/_596_ ( .A(\mlsu/_182_ ), .Z(\mem_rdata[30] ) );
BUF_X1 \mlsu/_597_ ( .A(\mlsu/_rdata[31] ), .Z(\mlsu/_023_ ) );
BUF_X1 \mlsu/_598_ ( .A(\mlsu/_183_ ), .Z(\mem_rdata[31] ) );
BUF_X1 \mlsu/_599_ ( .A(lsu_bready ), .Z(\mlsu/_071_ ) );
BUF_X1 \mlsu/_600_ ( .A(lsu_wvalid ), .Z(\mlsu/_107_ ) );
BUF_X1 \mlsu/_601_ ( .A(\mlsu/_030_ ), .Z(\mlsu/_237_ ) );
BUF_X1 \mlsu/_602_ ( .A(\mem_rdata[0] ), .Z(\mlsu/_159_ ) );
BUF_X1 \mlsu/_603_ ( .A(\lsu_rdata[0] ), .Z(\mlsu/_073_ ) );
BUF_X1 \mlsu/_604_ ( .A(\mlsu/_031_ ), .Z(\mlsu/_238_ ) );
BUF_X1 \mlsu/_605_ ( .A(\mem_rdata[1] ), .Z(\mlsu/_170_ ) );
BUF_X1 \mlsu/_606_ ( .A(\lsu_rdata[1] ), .Z(\mlsu/_084_ ) );
BUF_X1 \mlsu/_607_ ( .A(\mlsu/_032_ ), .Z(\mlsu/_239_ ) );
BUF_X1 \mlsu/_608_ ( .A(\mem_rdata[2] ), .Z(\mlsu/_181_ ) );
BUF_X1 \mlsu/_609_ ( .A(\lsu_rdata[2] ), .Z(\mlsu/_095_ ) );
BUF_X1 \mlsu/_610_ ( .A(\mlsu/_033_ ), .Z(\mlsu/_240_ ) );
BUF_X1 \mlsu/_611_ ( .A(\mem_rdata[3] ), .Z(\mlsu/_184_ ) );
BUF_X1 \mlsu/_612_ ( .A(\lsu_rdata[3] ), .Z(\mlsu/_098_ ) );
BUF_X1 \mlsu/_613_ ( .A(\mlsu/_034_ ), .Z(\mlsu/_241_ ) );
BUF_X1 \mlsu/_614_ ( .A(\mem_rdata[4] ), .Z(\mlsu/_185_ ) );
BUF_X1 \mlsu/_615_ ( .A(\lsu_rdata[4] ), .Z(\mlsu/_099_ ) );
BUF_X1 \mlsu/_616_ ( .A(\mlsu/_035_ ), .Z(\mlsu/_242_ ) );
BUF_X1 \mlsu/_617_ ( .A(\mem_rdata[5] ), .Z(\mlsu/_186_ ) );
BUF_X1 \mlsu/_618_ ( .A(\lsu_rdata[5] ), .Z(\mlsu/_100_ ) );
BUF_X1 \mlsu/_619_ ( .A(\mlsu/_036_ ), .Z(\mlsu/_243_ ) );
BUF_X1 \mlsu/_620_ ( .A(\mem_rdata[6] ), .Z(\mlsu/_187_ ) );
BUF_X1 \mlsu/_621_ ( .A(\lsu_rdata[6] ), .Z(\mlsu/_101_ ) );
BUF_X1 \mlsu/_622_ ( .A(\mlsu/_037_ ), .Z(\mlsu/_244_ ) );
BUF_X1 \mlsu/_623_ ( .A(\lsu_rdata[7] ), .Z(\mlsu/_102_ ) );
BUF_X1 \mlsu/_624_ ( .A(\mlsu/_038_ ), .Z(\mlsu/_245_ ) );
BUF_X1 \mlsu/_625_ ( .A(\lsu_rdata[8] ), .Z(\mlsu/_103_ ) );
BUF_X1 \mlsu/_626_ ( .A(\mlsu/_039_ ), .Z(\mlsu/_246_ ) );
BUF_X1 \mlsu/_627_ ( .A(\lsu_rdata[9] ), .Z(\mlsu/_104_ ) );
BUF_X1 \mlsu/_628_ ( .A(\mlsu/_040_ ), .Z(\mlsu/_247_ ) );
BUF_X1 \mlsu/_629_ ( .A(\lsu_rdata[10] ), .Z(\mlsu/_074_ ) );
BUF_X1 \mlsu/_630_ ( .A(\mlsu/_041_ ), .Z(\mlsu/_248_ ) );
BUF_X1 \mlsu/_631_ ( .A(\lsu_rdata[11] ), .Z(\mlsu/_075_ ) );
BUF_X1 \mlsu/_632_ ( .A(\mlsu/_042_ ), .Z(\mlsu/_249_ ) );
BUF_X1 \mlsu/_633_ ( .A(\lsu_rdata[12] ), .Z(\mlsu/_076_ ) );
BUF_X1 \mlsu/_634_ ( .A(\mlsu/_043_ ), .Z(\mlsu/_250_ ) );
BUF_X1 \mlsu/_635_ ( .A(\lsu_rdata[13] ), .Z(\mlsu/_077_ ) );
BUF_X1 \mlsu/_636_ ( .A(\mlsu/_044_ ), .Z(\mlsu/_251_ ) );
BUF_X1 \mlsu/_637_ ( .A(\lsu_rdata[14] ), .Z(\mlsu/_078_ ) );
BUF_X1 \mlsu/_638_ ( .A(\mlsu/_045_ ), .Z(\mlsu/_252_ ) );
BUF_X1 \mlsu/_639_ ( .A(\lsu_rdata[15] ), .Z(\mlsu/_079_ ) );
BUF_X1 \mlsu/_640_ ( .A(\mlsu/_046_ ), .Z(\mlsu/_253_ ) );
BUF_X1 \mlsu/_641_ ( .A(\lsu_rdata[16] ), .Z(\mlsu/_080_ ) );
BUF_X1 \mlsu/_642_ ( .A(\mlsu/_047_ ), .Z(\mlsu/_254_ ) );
BUF_X1 \mlsu/_643_ ( .A(\lsu_rdata[17] ), .Z(\mlsu/_081_ ) );
BUF_X1 \mlsu/_644_ ( .A(\mlsu/_048_ ), .Z(\mlsu/_255_ ) );
BUF_X1 \mlsu/_645_ ( .A(\lsu_rdata[18] ), .Z(\mlsu/_082_ ) );
BUF_X1 \mlsu/_646_ ( .A(\mlsu/_049_ ), .Z(\mlsu/_256_ ) );
BUF_X1 \mlsu/_647_ ( .A(\lsu_rdata[19] ), .Z(\mlsu/_083_ ) );
BUF_X1 \mlsu/_648_ ( .A(\mlsu/_050_ ), .Z(\mlsu/_257_ ) );
BUF_X1 \mlsu/_649_ ( .A(\lsu_rdata[20] ), .Z(\mlsu/_085_ ) );
BUF_X1 \mlsu/_650_ ( .A(\mlsu/_051_ ), .Z(\mlsu/_258_ ) );
BUF_X1 \mlsu/_651_ ( .A(\lsu_rdata[21] ), .Z(\mlsu/_086_ ) );
BUF_X1 \mlsu/_652_ ( .A(\mlsu/_052_ ), .Z(\mlsu/_259_ ) );
BUF_X1 \mlsu/_653_ ( .A(\lsu_rdata[22] ), .Z(\mlsu/_087_ ) );
BUF_X1 \mlsu/_654_ ( .A(\mlsu/_053_ ), .Z(\mlsu/_260_ ) );
BUF_X1 \mlsu/_655_ ( .A(\lsu_rdata[23] ), .Z(\mlsu/_088_ ) );
BUF_X1 \mlsu/_656_ ( .A(\mlsu/_054_ ), .Z(\mlsu/_261_ ) );
BUF_X1 \mlsu/_657_ ( .A(\lsu_rdata[24] ), .Z(\mlsu/_089_ ) );
BUF_X1 \mlsu/_658_ ( .A(\mlsu/_055_ ), .Z(\mlsu/_262_ ) );
BUF_X1 \mlsu/_659_ ( .A(\lsu_rdata[25] ), .Z(\mlsu/_090_ ) );
BUF_X1 \mlsu/_660_ ( .A(\mlsu/_056_ ), .Z(\mlsu/_263_ ) );
BUF_X1 \mlsu/_661_ ( .A(\lsu_rdata[26] ), .Z(\mlsu/_091_ ) );
BUF_X1 \mlsu/_662_ ( .A(\mlsu/_057_ ), .Z(\mlsu/_264_ ) );
BUF_X1 \mlsu/_663_ ( .A(\lsu_rdata[27] ), .Z(\mlsu/_092_ ) );
BUF_X1 \mlsu/_664_ ( .A(\mlsu/_058_ ), .Z(\mlsu/_265_ ) );
BUF_X1 \mlsu/_665_ ( .A(\lsu_rdata[28] ), .Z(\mlsu/_093_ ) );
BUF_X1 \mlsu/_666_ ( .A(\mlsu/_059_ ), .Z(\mlsu/_266_ ) );
BUF_X1 \mlsu/_667_ ( .A(\lsu_rdata[29] ), .Z(\mlsu/_094_ ) );
BUF_X1 \mlsu/_668_ ( .A(\mlsu/_060_ ), .Z(\mlsu/_267_ ) );
BUF_X1 \mlsu/_669_ ( .A(\lsu_rdata[30] ), .Z(\mlsu/_096_ ) );
BUF_X1 \mlsu/_670_ ( .A(\mlsu/_061_ ), .Z(\mlsu/_268_ ) );
BUF_X1 \mlsu/_671_ ( .A(\lsu_rdata[31] ), .Z(\mlsu/_097_ ) );
BUF_X1 \mlsu/_672_ ( .A(\mlsu/_062_ ), .Z(\mlsu/_269_ ) );
BUF_X1 \mlsu/_673_ ( .A(\mlsu/_026_ ), .Z(\mlsu/_233_ ) );
BUF_X1 \mlsu/_674_ ( .A(\mlsu/_027_ ), .Z(\mlsu/_234_ ) );
BUF_X1 \mlsu/_675_ ( .A(\mlsu/_028_ ), .Z(\mlsu/_235_ ) );
BUF_X1 \mlsu/_676_ ( .A(\mlsu/_029_ ), .Z(\mlsu/_236_ ) );
AND2_X2 \mpc/_327_ ( .A1(\mpc/_034_ ), .A2(\mpc/_263_ ), .ZN(\mpc/_035_ ) );
MUX2_X1 \mpc/_328_ ( .A(\mpc/_198_ ), .B(\mpc/_231_ ), .S(\mpc/_035_ ), .Z(\mpc/_036_ ) );
INV_X1 \mpc/_329_ ( .A(\mpc/_230_ ), .ZN(\mpc/_037_ ) );
AND2_X1 \mpc/_330_ ( .A1(\mpc/_036_ ), .A2(\mpc/_037_ ), .ZN(\mpc/_002_ ) );
MUX2_X1 \mpc/_331_ ( .A(\mpc/_209_ ), .B(\mpc/_242_ ), .S(\mpc/_035_ ), .Z(\mpc/_038_ ) );
AND2_X1 \mpc/_332_ ( .A1(\mpc/_038_ ), .A2(\mpc/_037_ ), .ZN(\mpc/_003_ ) );
INV_X1 \mpc/_333_ ( .A(\mpc/_263_ ), .ZN(\mpc/_039_ ) );
BUF_X4 \mpc/_334_ ( .A(\mpc/_039_ ), .Z(\mpc/_040_ ) );
AOI22_X1 \mpc/_335_ ( .A1(\mpc/_035_ ), .A2(\mpc/_253_ ), .B1(\mpc/_040_ ), .B2(\mpc/_220_ ), .ZN(\mpc/_041_ ) );
INV_X1 \mpc/_336_ ( .A(\mpc/_034_ ), .ZN(\mpc/_042_ ) );
NAND3_X1 \mpc/_337_ ( .A1(\mpc/_042_ ), .A2(\mpc/_263_ ), .A3(\mpc/_001_ ), .ZN(\mpc/_043_ ) );
AOI21_X1 \mpc/_338_ ( .A(\mpc/_230_ ), .B1(\mpc/_041_ ), .B2(\mpc/_043_ ), .ZN(\mpc/_004_ ) );
AND2_X4 \mpc/_339_ ( .A1(\mpc/_223_ ), .A2(\mpc/_220_ ), .ZN(\mpc/_044_ ) );
NOR2_X1 \mpc/_340_ ( .A1(\mpc/_223_ ), .A2(\mpc/_220_ ), .ZN(\mpc/_045_ ) );
OAI21_X1 \mpc/_341_ ( .A(\mpc/_042_ ), .B1(\mpc/_044_ ), .B2(\mpc/_045_ ), .ZN(\mpc/_046_ ) );
OAI211_X2 \mpc/_342_ ( .A(\mpc/_046_ ), .B(\mpc/_263_ ), .C1(\mpc/_042_ ), .C2(\mpc/_256_ ), .ZN(\mpc/_047_ ) );
NAND2_X1 \mpc/_343_ ( .A1(\mpc/_040_ ), .A2(\mpc/_223_ ), .ZN(\mpc/_048_ ) );
AOI21_X1 \mpc/_344_ ( .A(\mpc/_230_ ), .B1(\mpc/_047_ ), .B2(\mpc/_048_ ), .ZN(\mpc/_005_ ) );
NAND2_X1 \mpc/_345_ ( .A1(\mpc/_040_ ), .A2(\mpc/_224_ ), .ZN(\mpc/_049_ ) );
AND2_X4 \mpc/_346_ ( .A1(\mpc/_044_ ), .A2(\mpc/_224_ ), .ZN(\mpc/_050_ ) );
NOR2_X1 \mpc/_347_ ( .A1(\mpc/_039_ ), .A2(\mpc/_034_ ), .ZN(\mpc/_051_ ) );
INV_X1 \mpc/_348_ ( .A(\mpc/_051_ ), .ZN(\mpc/_052_ ) );
BUF_X4 \mpc/_349_ ( .A(\mpc/_052_ ), .Z(\mpc/_053_ ) );
OAI21_X1 \mpc/_350_ ( .A(\mpc/_049_ ), .B1(\mpc/_050_ ), .B2(\mpc/_053_ ), .ZN(\mpc/_054_ ) );
OAI21_X1 \mpc/_351_ ( .A(\mpc/_054_ ), .B1(\mpc/_224_ ), .B2(\mpc/_044_ ), .ZN(\mpc/_055_ ) );
NAND3_X1 \mpc/_352_ ( .A1(\mpc/_034_ ), .A2(\mpc/_263_ ), .A3(\mpc/_257_ ), .ZN(\mpc/_056_ ) );
AOI21_X1 \mpc/_353_ ( .A(\mpc/_230_ ), .B1(\mpc/_055_ ), .B2(\mpc/_056_ ), .ZN(\mpc/_006_ ) );
NAND2_X1 \mpc/_354_ ( .A1(\mpc/_040_ ), .A2(\mpc/_225_ ), .ZN(\mpc/_057_ ) );
AND2_X4 \mpc/_355_ ( .A1(\mpc/_050_ ), .A2(\mpc/_225_ ), .ZN(\mpc/_058_ ) );
OAI21_X1 \mpc/_356_ ( .A(\mpc/_057_ ), .B1(\mpc/_058_ ), .B2(\mpc/_053_ ), .ZN(\mpc/_059_ ) );
OAI21_X1 \mpc/_357_ ( .A(\mpc/_059_ ), .B1(\mpc/_225_ ), .B2(\mpc/_050_ ), .ZN(\mpc/_060_ ) );
NAND3_X1 \mpc/_358_ ( .A1(\mpc/_034_ ), .A2(\mpc/_263_ ), .A3(\mpc/_258_ ), .ZN(\mpc/_061_ ) );
AOI21_X1 \mpc/_359_ ( .A(\mpc/_230_ ), .B1(\mpc/_060_ ), .B2(\mpc/_061_ ), .ZN(\mpc/_007_ ) );
NAND2_X1 \mpc/_360_ ( .A1(\mpc/_040_ ), .A2(\mpc/_226_ ), .ZN(\mpc/_062_ ) );
AND2_X4 \mpc/_361_ ( .A1(\mpc/_058_ ), .A2(\mpc/_226_ ), .ZN(\mpc/_063_ ) );
OAI21_X1 \mpc/_362_ ( .A(\mpc/_062_ ), .B1(\mpc/_063_ ), .B2(\mpc/_053_ ), .ZN(\mpc/_064_ ) );
OAI21_X1 \mpc/_363_ ( .A(\mpc/_064_ ), .B1(\mpc/_226_ ), .B2(\mpc/_058_ ), .ZN(\mpc/_065_ ) );
NAND3_X1 \mpc/_364_ ( .A1(\mpc/_034_ ), .A2(\mpc/_263_ ), .A3(\mpc/_259_ ), .ZN(\mpc/_066_ ) );
AOI21_X1 \mpc/_365_ ( .A(\mpc/_230_ ), .B1(\mpc/_065_ ), .B2(\mpc/_066_ ), .ZN(\mpc/_008_ ) );
NAND2_X1 \mpc/_366_ ( .A1(\mpc/_040_ ), .A2(\mpc/_227_ ), .ZN(\mpc/_067_ ) );
AND2_X4 \mpc/_367_ ( .A1(\mpc/_063_ ), .A2(\mpc/_227_ ), .ZN(\mpc/_068_ ) );
OAI21_X1 \mpc/_368_ ( .A(\mpc/_067_ ), .B1(\mpc/_068_ ), .B2(\mpc/_053_ ), .ZN(\mpc/_069_ ) );
OAI21_X1 \mpc/_369_ ( .A(\mpc/_069_ ), .B1(\mpc/_227_ ), .B2(\mpc/_063_ ), .ZN(\mpc/_070_ ) );
NAND3_X1 \mpc/_370_ ( .A1(\mpc/_034_ ), .A2(\mpc/_263_ ), .A3(\mpc/_260_ ), .ZN(\mpc/_071_ ) );
AOI21_X1 \mpc/_371_ ( .A(\mpc/_230_ ), .B1(\mpc/_070_ ), .B2(\mpc/_071_ ), .ZN(\mpc/_009_ ) );
BUF_X2 \mpc/_372_ ( .A(\mpc/_039_ ), .Z(\mpc/_072_ ) );
BUF_X4 \mpc/_373_ ( .A(\mpc/_072_ ), .Z(\mpc/_073_ ) );
NAND2_X1 \mpc/_374_ ( .A1(\mpc/_073_ ), .A2(\mpc/_228_ ), .ZN(\mpc/_074_ ) );
AND2_X4 \mpc/_375_ ( .A1(\mpc/_068_ ), .A2(\mpc/_228_ ), .ZN(\mpc/_075_ ) );
OAI21_X1 \mpc/_376_ ( .A(\mpc/_074_ ), .B1(\mpc/_075_ ), .B2(\mpc/_053_ ), .ZN(\mpc/_076_ ) );
OAI21_X1 \mpc/_377_ ( .A(\mpc/_076_ ), .B1(\mpc/_228_ ), .B2(\mpc/_068_ ), .ZN(\mpc/_077_ ) );
NAND3_X1 \mpc/_378_ ( .A1(\mpc/_034_ ), .A2(\mpc/_263_ ), .A3(\mpc/_261_ ), .ZN(\mpc/_078_ ) );
AOI21_X1 \mpc/_379_ ( .A(\mpc/_230_ ), .B1(\mpc/_077_ ), .B2(\mpc/_078_ ), .ZN(\mpc/_010_ ) );
BUF_X4 \mpc/_380_ ( .A(\mpc/_052_ ), .Z(\mpc/_079_ ) );
AOI21_X1 \mpc/_381_ ( .A(\mpc/_079_ ), .B1(\mpc/_075_ ), .B2(\mpc/_229_ ), .ZN(\mpc/_080_ ) );
AND2_X1 \mpc/_382_ ( .A1(\mpc/_072_ ), .A2(\mpc/_229_ ), .ZN(\mpc/_081_ ) );
OAI22_X1 \mpc/_383_ ( .A1(\mpc/_080_ ), .A2(\mpc/_081_ ), .B1(\mpc/_229_ ), .B2(\mpc/_075_ ), .ZN(\mpc/_082_ ) );
NAND3_X1 \mpc/_384_ ( .A1(\mpc/_034_ ), .A2(\mpc/_263_ ), .A3(\mpc/_262_ ), .ZN(\mpc/_083_ ) );
AOI21_X1 \mpc/_385_ ( .A(\mpc/_230_ ), .B1(\mpc/_082_ ), .B2(\mpc/_083_ ), .ZN(\mpc/_011_ ) );
NAND2_X1 \mpc/_386_ ( .A1(\mpc/_073_ ), .A2(\mpc/_199_ ), .ZN(\mpc/_084_ ) );
AND2_X4 \mpc/_387_ ( .A1(\mpc/_075_ ), .A2(\mpc/_229_ ), .ZN(\mpc/_085_ ) );
AND2_X4 \mpc/_388_ ( .A1(\mpc/_085_ ), .A2(\mpc/_199_ ), .ZN(\mpc/_086_ ) );
OAI21_X1 \mpc/_389_ ( .A(\mpc/_084_ ), .B1(\mpc/_086_ ), .B2(\mpc/_053_ ), .ZN(\mpc/_087_ ) );
OAI21_X1 \mpc/_390_ ( .A(\mpc/_087_ ), .B1(\mpc/_199_ ), .B2(\mpc/_085_ ), .ZN(\mpc/_088_ ) );
NAND3_X1 \mpc/_391_ ( .A1(\mpc/_034_ ), .A2(\mpc/_263_ ), .A3(\mpc/_232_ ), .ZN(\mpc/_089_ ) );
AOI21_X1 \mpc/_392_ ( .A(\mpc/_230_ ), .B1(\mpc/_088_ ), .B2(\mpc/_089_ ), .ZN(\mpc/_012_ ) );
NAND2_X1 \mpc/_393_ ( .A1(\mpc/_073_ ), .A2(\mpc/_200_ ), .ZN(\mpc/_090_ ) );
AND2_X4 \mpc/_394_ ( .A1(\mpc/_086_ ), .A2(\mpc/_200_ ), .ZN(\mpc/_091_ ) );
OAI21_X1 \mpc/_395_ ( .A(\mpc/_090_ ), .B1(\mpc/_091_ ), .B2(\mpc/_053_ ), .ZN(\mpc/_092_ ) );
OAI21_X1 \mpc/_396_ ( .A(\mpc/_092_ ), .B1(\mpc/_200_ ), .B2(\mpc/_086_ ), .ZN(\mpc/_093_ ) );
NAND3_X1 \mpc/_397_ ( .A1(\mpc/_034_ ), .A2(\mpc/_263_ ), .A3(\mpc/_233_ ), .ZN(\mpc/_094_ ) );
AOI21_X1 \mpc/_398_ ( .A(\mpc/_230_ ), .B1(\mpc/_093_ ), .B2(\mpc/_094_ ), .ZN(\mpc/_013_ ) );
NAND2_X1 \mpc/_399_ ( .A1(\mpc/_073_ ), .A2(\mpc/_201_ ), .ZN(\mpc/_095_ ) );
AND2_X4 \mpc/_400_ ( .A1(\mpc/_091_ ), .A2(\mpc/_201_ ), .ZN(\mpc/_096_ ) );
OAI21_X1 \mpc/_401_ ( .A(\mpc/_095_ ), .B1(\mpc/_096_ ), .B2(\mpc/_053_ ), .ZN(\mpc/_097_ ) );
OAI21_X1 \mpc/_402_ ( .A(\mpc/_097_ ), .B1(\mpc/_201_ ), .B2(\mpc/_091_ ), .ZN(\mpc/_098_ ) );
NAND3_X1 \mpc/_403_ ( .A1(\mpc/_034_ ), .A2(\mpc/_263_ ), .A3(\mpc/_234_ ), .ZN(\mpc/_099_ ) );
AOI21_X1 \mpc/_404_ ( .A(\mpc/_230_ ), .B1(\mpc/_098_ ), .B2(\mpc/_099_ ), .ZN(\mpc/_014_ ) );
AOI21_X1 \mpc/_405_ ( .A(\mpc/_052_ ), .B1(\mpc/_096_ ), .B2(\mpc/_202_ ), .ZN(\mpc/_100_ ) );
AND2_X1 \mpc/_406_ ( .A1(\mpc/_072_ ), .A2(\mpc/_202_ ), .ZN(\mpc/_101_ ) );
OAI22_X1 \mpc/_407_ ( .A1(\mpc/_100_ ), .A2(\mpc/_101_ ), .B1(\mpc/_202_ ), .B2(\mpc/_096_ ), .ZN(\mpc/_102_ ) );
NAND3_X1 \mpc/_408_ ( .A1(\mpc/_034_ ), .A2(\mpc/_263_ ), .A3(\mpc/_235_ ), .ZN(\mpc/_103_ ) );
AOI21_X1 \mpc/_409_ ( .A(\mpc/_230_ ), .B1(\mpc/_102_ ), .B2(\mpc/_103_ ), .ZN(\mpc/_015_ ) );
NAND2_X1 \mpc/_410_ ( .A1(\mpc/_073_ ), .A2(\mpc/_203_ ), .ZN(\mpc/_104_ ) );
AND2_X4 \mpc/_411_ ( .A1(\mpc/_096_ ), .A2(\mpc/_202_ ), .ZN(\mpc/_105_ ) );
AND2_X1 \mpc/_412_ ( .A1(\mpc/_105_ ), .A2(\mpc/_203_ ), .ZN(\mpc/_106_ ) );
OAI21_X1 \mpc/_413_ ( .A(\mpc/_104_ ), .B1(\mpc/_106_ ), .B2(\mpc/_053_ ), .ZN(\mpc/_107_ ) );
OAI21_X1 \mpc/_414_ ( .A(\mpc/_107_ ), .B1(\mpc/_203_ ), .B2(\mpc/_105_ ), .ZN(\mpc/_108_ ) );
NAND3_X1 \mpc/_415_ ( .A1(\mpc/_034_ ), .A2(\mpc/_263_ ), .A3(\mpc/_236_ ), .ZN(\mpc/_109_ ) );
AOI21_X1 \mpc/_416_ ( .A(\mpc/_230_ ), .B1(\mpc/_108_ ), .B2(\mpc/_109_ ), .ZN(\mpc/_016_ ) );
NAND2_X1 \mpc/_417_ ( .A1(\mpc/_073_ ), .A2(\mpc/_204_ ), .ZN(\mpc/_110_ ) );
AND2_X1 \mpc/_418_ ( .A1(\mpc/_203_ ), .A2(\mpc/_204_ ), .ZN(\mpc/_111_ ) );
AND2_X1 \mpc/_419_ ( .A1(\mpc/_105_ ), .A2(\mpc/_111_ ), .ZN(\mpc/_112_ ) );
OAI21_X1 \mpc/_420_ ( .A(\mpc/_110_ ), .B1(\mpc/_112_ ), .B2(\mpc/_079_ ), .ZN(\mpc/_113_ ) );
OAI21_X1 \mpc/_421_ ( .A(\mpc/_113_ ), .B1(\mpc/_204_ ), .B2(\mpc/_106_ ), .ZN(\mpc/_114_ ) );
NAND3_X1 \mpc/_422_ ( .A1(\mpc/_034_ ), .A2(\mpc/_263_ ), .A3(\mpc/_237_ ), .ZN(\mpc/_115_ ) );
AOI21_X1 \mpc/_423_ ( .A(\mpc/_230_ ), .B1(\mpc/_114_ ), .B2(\mpc/_115_ ), .ZN(\mpc/_017_ ) );
AND2_X1 \mpc/_424_ ( .A1(\mpc/_112_ ), .A2(\mpc/_205_ ), .ZN(\mpc/_116_ ) );
INV_X1 \mpc/_425_ ( .A(\mpc/_205_ ), .ZN(\mpc/_117_ ) );
OAI22_X1 \mpc/_426_ ( .A1(\mpc/_116_ ), .A2(\mpc/_079_ ), .B1(\mpc/_263_ ), .B2(\mpc/_117_ ), .ZN(\mpc/_118_ ) );
AND3_X4 \mpc/_427_ ( .A1(\mpc/_105_ ), .A2(\mpc/_203_ ), .A3(\mpc/_204_ ), .ZN(\mpc/_119_ ) );
OAI21_X1 \mpc/_428_ ( .A(\mpc/_118_ ), .B1(\mpc/_205_ ), .B2(\mpc/_119_ ), .ZN(\mpc/_120_ ) );
NAND3_X1 \mpc/_429_ ( .A1(\mpc/_034_ ), .A2(\mpc/_263_ ), .A3(\mpc/_238_ ), .ZN(\mpc/_121_ ) );
AOI21_X1 \mpc/_430_ ( .A(\mpc/_230_ ), .B1(\mpc/_120_ ), .B2(\mpc/_121_ ), .ZN(\mpc/_018_ ) );
AND2_X4 \mpc/_431_ ( .A1(\mpc/_119_ ), .A2(\mpc/_205_ ), .ZN(\mpc/_122_ ) );
AOI21_X1 \mpc/_432_ ( .A(\mpc/_052_ ), .B1(\mpc/_122_ ), .B2(\mpc/_206_ ), .ZN(\mpc/_123_ ) );
AND2_X1 \mpc/_433_ ( .A1(\mpc/_072_ ), .A2(\mpc/_206_ ), .ZN(\mpc/_124_ ) );
OAI22_X1 \mpc/_434_ ( .A1(\mpc/_123_ ), .A2(\mpc/_124_ ), .B1(\mpc/_206_ ), .B2(\mpc/_122_ ), .ZN(\mpc/_125_ ) );
NAND3_X1 \mpc/_435_ ( .A1(\mpc/_034_ ), .A2(\mpc/_263_ ), .A3(\mpc/_239_ ), .ZN(\mpc/_126_ ) );
AOI21_X1 \mpc/_436_ ( .A(\mpc/_230_ ), .B1(\mpc/_125_ ), .B2(\mpc/_126_ ), .ZN(\mpc/_019_ ) );
NAND2_X1 \mpc/_437_ ( .A1(\mpc/_073_ ), .A2(\mpc/_207_ ), .ZN(\mpc/_127_ ) );
AND2_X4 \mpc/_438_ ( .A1(\mpc/_122_ ), .A2(\mpc/_206_ ), .ZN(\mpc/_128_ ) );
AND2_X1 \mpc/_439_ ( .A1(\mpc/_128_ ), .A2(\mpc/_207_ ), .ZN(\mpc/_129_ ) );
OAI21_X1 \mpc/_440_ ( .A(\mpc/_127_ ), .B1(\mpc/_129_ ), .B2(\mpc/_079_ ), .ZN(\mpc/_130_ ) );
OAI21_X1 \mpc/_441_ ( .A(\mpc/_130_ ), .B1(\mpc/_207_ ), .B2(\mpc/_128_ ), .ZN(\mpc/_131_ ) );
NAND3_X1 \mpc/_442_ ( .A1(\mpc/_034_ ), .A2(\mpc/_263_ ), .A3(\mpc/_240_ ), .ZN(\mpc/_132_ ) );
AOI21_X1 \mpc/_443_ ( .A(\mpc/_230_ ), .B1(\mpc/_131_ ), .B2(\mpc/_132_ ), .ZN(\mpc/_020_ ) );
NAND2_X1 \mpc/_444_ ( .A1(\mpc/_073_ ), .A2(\mpc/_208_ ), .ZN(\mpc/_133_ ) );
AND2_X1 \mpc/_445_ ( .A1(\mpc/_207_ ), .A2(\mpc/_208_ ), .ZN(\mpc/_134_ ) );
AND2_X1 \mpc/_446_ ( .A1(\mpc/_128_ ), .A2(\mpc/_134_ ), .ZN(\mpc/_135_ ) );
OAI21_X1 \mpc/_447_ ( .A(\mpc/_133_ ), .B1(\mpc/_135_ ), .B2(\mpc/_079_ ), .ZN(\mpc/_136_ ) );
OAI21_X1 \mpc/_448_ ( .A(\mpc/_136_ ), .B1(\mpc/_208_ ), .B2(\mpc/_129_ ), .ZN(\mpc/_137_ ) );
NAND3_X1 \mpc/_449_ ( .A1(\mpc/_034_ ), .A2(\mpc/_263_ ), .A3(\mpc/_241_ ), .ZN(\mpc/_138_ ) );
AOI21_X1 \mpc/_450_ ( .A(\mpc/_230_ ), .B1(\mpc/_137_ ), .B2(\mpc/_138_ ), .ZN(\mpc/_021_ ) );
AOI21_X1 \mpc/_451_ ( .A(\mpc/_052_ ), .B1(\mpc/_135_ ), .B2(\mpc/_210_ ), .ZN(\mpc/_139_ ) );
AND2_X1 \mpc/_452_ ( .A1(\mpc/_072_ ), .A2(\mpc/_210_ ), .ZN(\mpc/_140_ ) );
AND3_X1 \mpc/_453_ ( .A1(\mpc/_128_ ), .A2(\mpc/_207_ ), .A3(\mpc/_208_ ), .ZN(\mpc/_141_ ) );
OAI22_X1 \mpc/_454_ ( .A1(\mpc/_139_ ), .A2(\mpc/_140_ ), .B1(\mpc/_210_ ), .B2(\mpc/_141_ ), .ZN(\mpc/_142_ ) );
NAND3_X1 \mpc/_455_ ( .A1(\mpc/_034_ ), .A2(\mpc/_263_ ), .A3(\mpc/_243_ ), .ZN(\mpc/_143_ ) );
AOI21_X1 \mpc/_456_ ( .A(\mpc/_230_ ), .B1(\mpc/_142_ ), .B2(\mpc/_143_ ), .ZN(\mpc/_022_ ) );
AND2_X1 \mpc/_457_ ( .A1(\mpc/_135_ ), .A2(\mpc/_210_ ), .ZN(\mpc/_144_ ) );
AND2_X1 \mpc/_458_ ( .A1(\mpc/_072_ ), .A2(\mpc/_211_ ), .ZN(\mpc/_145_ ) );
AND3_X1 \mpc/_459_ ( .A1(\mpc/_134_ ), .A2(\mpc/_210_ ), .A3(\mpc/_211_ ), .ZN(\mpc/_146_ ) );
AOI21_X1 \mpc/_460_ ( .A(\mpc/_052_ ), .B1(\mpc/_128_ ), .B2(\mpc/_146_ ), .ZN(\mpc/_147_ ) );
OAI22_X1 \mpc/_461_ ( .A1(\mpc/_144_ ), .A2(\mpc/_211_ ), .B1(\mpc/_145_ ), .B2(\mpc/_147_ ), .ZN(\mpc/_148_ ) );
NAND3_X1 \mpc/_462_ ( .A1(\mpc/_034_ ), .A2(\mpc/_263_ ), .A3(\mpc/_244_ ), .ZN(\mpc/_149_ ) );
AOI21_X1 \mpc/_463_ ( .A(\mpc/_230_ ), .B1(\mpc/_148_ ), .B2(\mpc/_149_ ), .ZN(\mpc/_023_ ) );
NAND2_X1 \mpc/_464_ ( .A1(\mpc/_073_ ), .A2(\mpc/_212_ ), .ZN(\mpc/_150_ ) );
AND2_X1 \mpc/_465_ ( .A1(\mpc/_128_ ), .A2(\mpc/_146_ ), .ZN(\mpc/_151_ ) );
AND2_X1 \mpc/_466_ ( .A1(\mpc/_151_ ), .A2(\mpc/_212_ ), .ZN(\mpc/_152_ ) );
OAI21_X1 \mpc/_467_ ( .A(\mpc/_150_ ), .B1(\mpc/_152_ ), .B2(\mpc/_079_ ), .ZN(\mpc/_153_ ) );
OAI21_X1 \mpc/_468_ ( .A(\mpc/_153_ ), .B1(\mpc/_212_ ), .B2(\mpc/_151_ ), .ZN(\mpc/_154_ ) );
NAND3_X1 \mpc/_469_ ( .A1(\mpc/_034_ ), .A2(\mpc/_263_ ), .A3(\mpc/_245_ ), .ZN(\mpc/_155_ ) );
AOI21_X1 \mpc/_470_ ( .A(\mpc/_230_ ), .B1(\mpc/_154_ ), .B2(\mpc/_155_ ), .ZN(\mpc/_024_ ) );
NAND2_X1 \mpc/_471_ ( .A1(\mpc/_073_ ), .A2(\mpc/_213_ ), .ZN(\mpc/_156_ ) );
AND2_X1 \mpc/_472_ ( .A1(\mpc/_212_ ), .A2(\mpc/_213_ ), .ZN(\mpc/_157_ ) );
AND2_X1 \mpc/_473_ ( .A1(\mpc/_151_ ), .A2(\mpc/_157_ ), .ZN(\mpc/_158_ ) );
OAI21_X1 \mpc/_474_ ( .A(\mpc/_156_ ), .B1(\mpc/_158_ ), .B2(\mpc/_079_ ), .ZN(\mpc/_159_ ) );
OAI21_X1 \mpc/_475_ ( .A(\mpc/_159_ ), .B1(\mpc/_213_ ), .B2(\mpc/_152_ ), .ZN(\mpc/_160_ ) );
NAND3_X1 \mpc/_476_ ( .A1(\mpc/_034_ ), .A2(\mpc/_263_ ), .A3(\mpc/_246_ ), .ZN(\mpc/_161_ ) );
AOI21_X1 \mpc/_477_ ( .A(\mpc/_230_ ), .B1(\mpc/_160_ ), .B2(\mpc/_161_ ), .ZN(\mpc/_025_ ) );
AOI21_X1 \mpc/_478_ ( .A(\mpc/_034_ ), .B1(\mpc/_158_ ), .B2(\mpc/_214_ ), .ZN(\mpc/_162_ ) );
OAI211_X2 \mpc/_479_ ( .A(\mpc/_162_ ), .B(\mpc/_263_ ), .C1(\mpc/_214_ ), .C2(\mpc/_158_ ), .ZN(\mpc/_163_ ) );
AOI22_X1 \mpc/_480_ ( .A1(\mpc/_035_ ), .A2(\mpc/_247_ ), .B1(\mpc/_040_ ), .B2(\mpc/_214_ ), .ZN(\mpc/_164_ ) );
AOI21_X1 \mpc/_481_ ( .A(\mpc/_230_ ), .B1(\mpc/_163_ ), .B2(\mpc/_164_ ), .ZN(\mpc/_026_ ) );
AND4_X1 \mpc/_482_ ( .A1(\mpc/_214_ ), .A2(\mpc/_146_ ), .A3(\mpc/_215_ ), .A4(\mpc/_157_ ), .ZN(\mpc/_165_ ) );
AND2_X4 \mpc/_483_ ( .A1(\mpc/_128_ ), .A2(\mpc/_165_ ), .ZN(\mpc/_166_ ) );
INV_X1 \mpc/_484_ ( .A(\mpc/_166_ ), .ZN(\mpc/_167_ ) );
AND2_X1 \mpc/_485_ ( .A1(\mpc/_158_ ), .A2(\mpc/_214_ ), .ZN(\mpc/_168_ ) );
OAI211_X2 \mpc/_486_ ( .A(\mpc/_051_ ), .B(\mpc/_167_ ), .C1(\mpc/_168_ ), .C2(\mpc/_215_ ), .ZN(\mpc/_169_ ) );
AOI22_X1 \mpc/_487_ ( .A1(\mpc/_035_ ), .A2(\mpc/_248_ ), .B1(\mpc/_040_ ), .B2(\mpc/_215_ ), .ZN(\mpc/_170_ ) );
AOI21_X1 \mpc/_488_ ( .A(\mpc/_230_ ), .B1(\mpc/_169_ ), .B2(\mpc/_170_ ), .ZN(\mpc/_027_ ) );
NAND2_X1 \mpc/_489_ ( .A1(\mpc/_072_ ), .A2(\mpc/_216_ ), .ZN(\mpc/_171_ ) );
AND2_X1 \mpc/_490_ ( .A1(\mpc/_166_ ), .A2(\mpc/_216_ ), .ZN(\mpc/_172_ ) );
OAI21_X1 \mpc/_491_ ( .A(\mpc/_171_ ), .B1(\mpc/_172_ ), .B2(\mpc/_079_ ), .ZN(\mpc/_173_ ) );
OAI21_X1 \mpc/_492_ ( .A(\mpc/_173_ ), .B1(\mpc/_216_ ), .B2(\mpc/_166_ ), .ZN(\mpc/_174_ ) );
NAND3_X1 \mpc/_493_ ( .A1(\mpc/_034_ ), .A2(\mpc/_263_ ), .A3(\mpc/_249_ ), .ZN(\mpc/_175_ ) );
AOI21_X1 \mpc/_494_ ( .A(\mpc/_230_ ), .B1(\mpc/_174_ ), .B2(\mpc/_175_ ), .ZN(\mpc/_028_ ) );
NAND2_X1 \mpc/_495_ ( .A1(\mpc/_072_ ), .A2(\mpc/_217_ ), .ZN(\mpc/_176_ ) );
AND2_X1 \mpc/_496_ ( .A1(\mpc/_216_ ), .A2(\mpc/_217_ ), .ZN(\mpc/_177_ ) );
AND2_X4 \mpc/_497_ ( .A1(\mpc/_166_ ), .A2(\mpc/_177_ ), .ZN(\mpc/_178_ ) );
OAI21_X1 \mpc/_498_ ( .A(\mpc/_176_ ), .B1(\mpc/_178_ ), .B2(\mpc/_079_ ), .ZN(\mpc/_179_ ) );
OAI21_X1 \mpc/_499_ ( .A(\mpc/_179_ ), .B1(\mpc/_217_ ), .B2(\mpc/_172_ ), .ZN(\mpc/_180_ ) );
NAND3_X1 \mpc/_500_ ( .A1(\mpc/_034_ ), .A2(\mpc/_263_ ), .A3(\mpc/_250_ ), .ZN(\mpc/_181_ ) );
AOI21_X1 \mpc/_501_ ( .A(\mpc/_230_ ), .B1(\mpc/_180_ ), .B2(\mpc/_181_ ), .ZN(\mpc/_029_ ) );
AOI21_X1 \mpc/_502_ ( .A(\mpc/_034_ ), .B1(\mpc/_178_ ), .B2(\mpc/_218_ ), .ZN(\mpc/_182_ ) );
OAI211_X2 \mpc/_503_ ( .A(\mpc/_182_ ), .B(\mpc/_263_ ), .C1(\mpc/_218_ ), .C2(\mpc/_178_ ), .ZN(\mpc/_183_ ) );
AOI22_X1 \mpc/_504_ ( .A1(\mpc/_035_ ), .A2(\mpc/_251_ ), .B1(\mpc/_040_ ), .B2(\mpc/_218_ ), .ZN(\mpc/_184_ ) );
AOI21_X1 \mpc/_505_ ( .A(\mpc/_230_ ), .B1(\mpc/_183_ ), .B2(\mpc/_184_ ), .ZN(\mpc/_030_ ) );
NAND2_X1 \mpc/_506_ ( .A1(\mpc/_072_ ), .A2(\mpc/_219_ ), .ZN(\mpc/_185_ ) );
AND3_X4 \mpc/_507_ ( .A1(\mpc/_178_ ), .A2(\mpc/_218_ ), .A3(\mpc/_219_ ), .ZN(\mpc/_186_ ) );
OAI21_X1 \mpc/_508_ ( .A(\mpc/_185_ ), .B1(\mpc/_186_ ), .B2(\mpc/_079_ ), .ZN(\mpc/_187_ ) );
AND2_X1 \mpc/_509_ ( .A1(\mpc/_178_ ), .A2(\mpc/_218_ ), .ZN(\mpc/_188_ ) );
OAI21_X1 \mpc/_510_ ( .A(\mpc/_187_ ), .B1(\mpc/_219_ ), .B2(\mpc/_188_ ), .ZN(\mpc/_189_ ) );
NAND3_X1 \mpc/_511_ ( .A1(\mpc/_034_ ), .A2(\mpc/_263_ ), .A3(\mpc/_252_ ), .ZN(\mpc/_190_ ) );
AOI21_X1 \mpc/_512_ ( .A(\mpc/_230_ ), .B1(\mpc/_189_ ), .B2(\mpc/_190_ ), .ZN(\mpc/_031_ ) );
AND2_X4 \mpc/_513_ ( .A1(\mpc/_186_ ), .A2(\mpc/_221_ ), .ZN(\mpc/_191_ ) );
INV_X1 \mpc/_514_ ( .A(\mpc/_191_ ), .ZN(\mpc/_192_ ) );
AND3_X1 \mpc/_515_ ( .A1(\mpc/_178_ ), .A2(\mpc/_218_ ), .A3(\mpc/_219_ ), .ZN(\mpc/_193_ ) );
OAI211_X2 \mpc/_516_ ( .A(\mpc/_192_ ), .B(\mpc/_051_ ), .C1(\mpc/_221_ ), .C2(\mpc/_193_ ), .ZN(\mpc/_194_ ) );
AOI22_X1 \mpc/_517_ ( .A1(\mpc/_035_ ), .A2(\mpc/_254_ ), .B1(\mpc/_040_ ), .B2(\mpc/_221_ ), .ZN(\mpc/_195_ ) );
AOI21_X1 \mpc/_518_ ( .A(\mpc/_230_ ), .B1(\mpc/_194_ ), .B2(\mpc/_195_ ), .ZN(\mpc/_032_ ) );
AOI221_X4 \mpc/_519_ ( .A(\mpc/_230_ ), .B1(\mpc/_072_ ), .B2(\mpc/_222_ ), .C1(\mpc/_035_ ), .C2(\mpc/_255_ ), .ZN(\mpc/_196_ ) );
XNOR2_X2 \mpc/_520_ ( .A(\mpc/_191_ ), .B(\mpc/_222_ ), .ZN(\mpc/_197_ ) );
OAI21_X1 \mpc/_521_ ( .A(\mpc/_196_ ), .B1(\mpc/_197_ ), .B2(\mpc/_053_ ), .ZN(\mpc/_033_ ) );
DFF_X1 \mpc/_522_ ( .CK(clk ), .D(\mpc/_295_ ), .Q(\pc[0] ), .QN(\mpc/_294_ ) );
DFF_X1 \mpc/_523_ ( .CK(clk ), .D(\mpc/_296_ ), .Q(\pc[1] ), .QN(\mpc/_293_ ) );
DFF_X1 \mpc/_524_ ( .CK(clk ), .D(\mpc/_297_ ), .Q(\pc[2] ), .QN(\mpc/_000_ ) );
DFF_X1 \mpc/_525_ ( .CK(clk ), .D(\mpc/_298_ ), .Q(\pc[3] ), .QN(\mpc/_292_ ) );
DFF_X1 \mpc/_526_ ( .CK(clk ), .D(\mpc/_299_ ), .Q(\pc[4] ), .QN(\mpc/_291_ ) );
DFF_X1 \mpc/_527_ ( .CK(clk ), .D(\mpc/_300_ ), .Q(\pc[5] ), .QN(\mpc/_290_ ) );
DFF_X1 \mpc/_528_ ( .CK(clk ), .D(\mpc/_301_ ), .Q(\pc[6] ), .QN(\mpc/_289_ ) );
DFF_X1 \mpc/_529_ ( .CK(clk ), .D(\mpc/_302_ ), .Q(\pc[7] ), .QN(\mpc/_288_ ) );
DFF_X1 \mpc/_530_ ( .CK(clk ), .D(\mpc/_303_ ), .Q(\pc[8] ), .QN(\mpc/_287_ ) );
DFF_X1 \mpc/_531_ ( .CK(clk ), .D(\mpc/_304_ ), .Q(\pc[9] ), .QN(\mpc/_286_ ) );
DFF_X1 \mpc/_532_ ( .CK(clk ), .D(\mpc/_305_ ), .Q(\pc[10] ), .QN(\mpc/_285_ ) );
DFF_X1 \mpc/_533_ ( .CK(clk ), .D(\mpc/_306_ ), .Q(\pc[11] ), .QN(\mpc/_284_ ) );
DFF_X1 \mpc/_534_ ( .CK(clk ), .D(\mpc/_307_ ), .Q(\pc[12] ), .QN(\mpc/_283_ ) );
DFF_X1 \mpc/_535_ ( .CK(clk ), .D(\mpc/_308_ ), .Q(\pc[13] ), .QN(\mpc/_282_ ) );
DFF_X1 \mpc/_536_ ( .CK(clk ), .D(\mpc/_309_ ), .Q(\pc[14] ), .QN(\mpc/_281_ ) );
DFF_X1 \mpc/_537_ ( .CK(clk ), .D(\mpc/_310_ ), .Q(\pc[15] ), .QN(\mpc/_280_ ) );
DFF_X1 \mpc/_538_ ( .CK(clk ), .D(\mpc/_311_ ), .Q(\pc[16] ), .QN(\mpc/_279_ ) );
DFF_X1 \mpc/_539_ ( .CK(clk ), .D(\mpc/_312_ ), .Q(\pc[17] ), .QN(\mpc/_278_ ) );
DFF_X1 \mpc/_540_ ( .CK(clk ), .D(\mpc/_313_ ), .Q(\pc[18] ), .QN(\mpc/_277_ ) );
DFF_X1 \mpc/_541_ ( .CK(clk ), .D(\mpc/_314_ ), .Q(\pc[19] ), .QN(\mpc/_276_ ) );
DFF_X1 \mpc/_542_ ( .CK(clk ), .D(\mpc/_315_ ), .Q(\pc[20] ), .QN(\mpc/_275_ ) );
DFF_X1 \mpc/_543_ ( .CK(clk ), .D(\mpc/_316_ ), .Q(\pc[21] ), .QN(\mpc/_274_ ) );
DFF_X1 \mpc/_544_ ( .CK(clk ), .D(\mpc/_317_ ), .Q(\pc[22] ), .QN(\mpc/_273_ ) );
DFF_X1 \mpc/_545_ ( .CK(clk ), .D(\mpc/_318_ ), .Q(\pc[23] ), .QN(\mpc/_272_ ) );
DFF_X1 \mpc/_546_ ( .CK(clk ), .D(\mpc/_319_ ), .Q(\pc[24] ), .QN(\mpc/_271_ ) );
DFF_X1 \mpc/_547_ ( .CK(clk ), .D(\mpc/_320_ ), .Q(\pc[25] ), .QN(\mpc/_270_ ) );
DFF_X1 \mpc/_548_ ( .CK(clk ), .D(\mpc/_321_ ), .Q(\pc[26] ), .QN(\mpc/_269_ ) );
DFF_X1 \mpc/_549_ ( .CK(clk ), .D(\mpc/_322_ ), .Q(\pc[27] ), .QN(\mpc/_268_ ) );
DFF_X1 \mpc/_550_ ( .CK(clk ), .D(\mpc/_323_ ), .Q(\pc[28] ), .QN(\mpc/_267_ ) );
DFF_X1 \mpc/_551_ ( .CK(clk ), .D(\mpc/_324_ ), .Q(\pc[29] ), .QN(\mpc/_266_ ) );
DFF_X1 \mpc/_552_ ( .CK(clk ), .D(\mpc/_325_ ), .Q(\pc[30] ), .QN(\mpc/_265_ ) );
DFF_X1 \mpc/_553_ ( .CK(clk ), .D(\mpc/_326_ ), .Q(\pc[31] ), .QN(\mpc/_264_ ) );
BUF_X1 \mpc/_554_ ( .A(jump ), .Z(\mpc/_034_ ) );
BUF_X1 \mpc/_555_ ( .A(pc_wen ), .Z(\mpc/_263_ ) );
BUF_X1 \mpc/_556_ ( .A(\upc[0] ), .Z(\mpc/_231_ ) );
BUF_X1 \mpc/_557_ ( .A(\upc[1] ), .Z(\mpc/_242_ ) );
BUF_X1 \mpc/_558_ ( .A(\mpc/_000_ ), .Z(\mpc/_001_ ) );
BUF_X1 \mpc/_559_ ( .A(\upc[2] ), .Z(\mpc/_253_ ) );
BUF_X1 \mpc/_560_ ( .A(\pc[3] ), .Z(\mpc/_223_ ) );
BUF_X1 \mpc/_561_ ( .A(\pc[2] ), .Z(\mpc/_220_ ) );
BUF_X1 \mpc/_562_ ( .A(\upc[3] ), .Z(\mpc/_256_ ) );
BUF_X1 \mpc/_563_ ( .A(\pc[4] ), .Z(\mpc/_224_ ) );
BUF_X1 \mpc/_564_ ( .A(\upc[4] ), .Z(\mpc/_257_ ) );
BUF_X1 \mpc/_565_ ( .A(\pc[5] ), .Z(\mpc/_225_ ) );
BUF_X1 \mpc/_566_ ( .A(\upc[5] ), .Z(\mpc/_258_ ) );
BUF_X1 \mpc/_567_ ( .A(\pc[6] ), .Z(\mpc/_226_ ) );
BUF_X1 \mpc/_568_ ( .A(\upc[6] ), .Z(\mpc/_259_ ) );
BUF_X1 \mpc/_569_ ( .A(\pc[7] ), .Z(\mpc/_227_ ) );
BUF_X1 \mpc/_570_ ( .A(\upc[7] ), .Z(\mpc/_260_ ) );
BUF_X1 \mpc/_571_ ( .A(\pc[8] ), .Z(\mpc/_228_ ) );
BUF_X1 \mpc/_572_ ( .A(\upc[8] ), .Z(\mpc/_261_ ) );
BUF_X1 \mpc/_573_ ( .A(\pc[9] ), .Z(\mpc/_229_ ) );
BUF_X1 \mpc/_574_ ( .A(\upc[9] ), .Z(\mpc/_262_ ) );
BUF_X1 \mpc/_575_ ( .A(\pc[10] ), .Z(\mpc/_199_ ) );
BUF_X1 \mpc/_576_ ( .A(\upc[10] ), .Z(\mpc/_232_ ) );
BUF_X1 \mpc/_577_ ( .A(\pc[11] ), .Z(\mpc/_200_ ) );
BUF_X1 \mpc/_578_ ( .A(\upc[11] ), .Z(\mpc/_233_ ) );
BUF_X1 \mpc/_579_ ( .A(\pc[12] ), .Z(\mpc/_201_ ) );
BUF_X1 \mpc/_580_ ( .A(\upc[12] ), .Z(\mpc/_234_ ) );
BUF_X1 \mpc/_581_ ( .A(\pc[13] ), .Z(\mpc/_202_ ) );
BUF_X1 \mpc/_582_ ( .A(\upc[13] ), .Z(\mpc/_235_ ) );
BUF_X1 \mpc/_583_ ( .A(\pc[14] ), .Z(\mpc/_203_ ) );
BUF_X1 \mpc/_584_ ( .A(\upc[14] ), .Z(\mpc/_236_ ) );
BUF_X1 \mpc/_585_ ( .A(\pc[15] ), .Z(\mpc/_204_ ) );
BUF_X1 \mpc/_586_ ( .A(\upc[15] ), .Z(\mpc/_237_ ) );
BUF_X1 \mpc/_587_ ( .A(\pc[16] ), .Z(\mpc/_205_ ) );
BUF_X1 \mpc/_588_ ( .A(\upc[16] ), .Z(\mpc/_238_ ) );
BUF_X1 \mpc/_589_ ( .A(\pc[17] ), .Z(\mpc/_206_ ) );
BUF_X1 \mpc/_590_ ( .A(\upc[17] ), .Z(\mpc/_239_ ) );
BUF_X1 \mpc/_591_ ( .A(\pc[18] ), .Z(\mpc/_207_ ) );
BUF_X1 \mpc/_592_ ( .A(\upc[18] ), .Z(\mpc/_240_ ) );
BUF_X1 \mpc/_593_ ( .A(\pc[19] ), .Z(\mpc/_208_ ) );
BUF_X1 \mpc/_594_ ( .A(\upc[19] ), .Z(\mpc/_241_ ) );
BUF_X1 \mpc/_595_ ( .A(\pc[20] ), .Z(\mpc/_210_ ) );
BUF_X1 \mpc/_596_ ( .A(\upc[20] ), .Z(\mpc/_243_ ) );
BUF_X1 \mpc/_597_ ( .A(\pc[21] ), .Z(\mpc/_211_ ) );
BUF_X1 \mpc/_598_ ( .A(\upc[21] ), .Z(\mpc/_244_ ) );
BUF_X1 \mpc/_599_ ( .A(\pc[22] ), .Z(\mpc/_212_ ) );
BUF_X1 \mpc/_600_ ( .A(\upc[22] ), .Z(\mpc/_245_ ) );
BUF_X1 \mpc/_601_ ( .A(\pc[23] ), .Z(\mpc/_213_ ) );
BUF_X1 \mpc/_602_ ( .A(\upc[23] ), .Z(\mpc/_246_ ) );
BUF_X1 \mpc/_603_ ( .A(\pc[24] ), .Z(\mpc/_214_ ) );
BUF_X1 \mpc/_604_ ( .A(\upc[24] ), .Z(\mpc/_247_ ) );
BUF_X1 \mpc/_605_ ( .A(\pc[25] ), .Z(\mpc/_215_ ) );
BUF_X1 \mpc/_606_ ( .A(\upc[25] ), .Z(\mpc/_248_ ) );
BUF_X1 \mpc/_607_ ( .A(\pc[26] ), .Z(\mpc/_216_ ) );
BUF_X1 \mpc/_608_ ( .A(\upc[26] ), .Z(\mpc/_249_ ) );
BUF_X1 \mpc/_609_ ( .A(\pc[27] ), .Z(\mpc/_217_ ) );
BUF_X1 \mpc/_610_ ( .A(\upc[27] ), .Z(\mpc/_250_ ) );
BUF_X1 \mpc/_611_ ( .A(\pc[28] ), .Z(\mpc/_218_ ) );
BUF_X1 \mpc/_612_ ( .A(\upc[28] ), .Z(\mpc/_251_ ) );
BUF_X1 \mpc/_613_ ( .A(\pc[29] ), .Z(\mpc/_219_ ) );
BUF_X1 \mpc/_614_ ( .A(\upc[29] ), .Z(\mpc/_252_ ) );
BUF_X1 \mpc/_615_ ( .A(\pc[30] ), .Z(\mpc/_221_ ) );
BUF_X1 \mpc/_616_ ( .A(\upc[30] ), .Z(\mpc/_254_ ) );
BUF_X1 \mpc/_617_ ( .A(\pc[31] ), .Z(\mpc/_222_ ) );
BUF_X1 \mpc/_618_ ( .A(\upc[31] ), .Z(\mpc/_255_ ) );
BUF_X1 \mpc/_619_ ( .A(\pc[0] ), .Z(\mpc/_198_ ) );
BUF_X1 \mpc/_620_ ( .A(\pc[1] ), .Z(\mpc/_209_ ) );
BUF_X1 \mpc/_621_ ( .A(rst ), .Z(\mpc/_230_ ) );
BUF_X1 \mpc/_622_ ( .A(\mpc/_002_ ), .Z(\mpc/_295_ ) );
BUF_X1 \mpc/_623_ ( .A(\mpc/_003_ ), .Z(\mpc/_296_ ) );
BUF_X1 \mpc/_624_ ( .A(\mpc/_004_ ), .Z(\mpc/_297_ ) );
BUF_X1 \mpc/_625_ ( .A(\mpc/_005_ ), .Z(\mpc/_298_ ) );
BUF_X1 \mpc/_626_ ( .A(\mpc/_006_ ), .Z(\mpc/_299_ ) );
BUF_X1 \mpc/_627_ ( .A(\mpc/_007_ ), .Z(\mpc/_300_ ) );
BUF_X1 \mpc/_628_ ( .A(\mpc/_008_ ), .Z(\mpc/_301_ ) );
BUF_X1 \mpc/_629_ ( .A(\mpc/_009_ ), .Z(\mpc/_302_ ) );
BUF_X1 \mpc/_630_ ( .A(\mpc/_010_ ), .Z(\mpc/_303_ ) );
BUF_X1 \mpc/_631_ ( .A(\mpc/_011_ ), .Z(\mpc/_304_ ) );
BUF_X1 \mpc/_632_ ( .A(\mpc/_012_ ), .Z(\mpc/_305_ ) );
BUF_X1 \mpc/_633_ ( .A(\mpc/_013_ ), .Z(\mpc/_306_ ) );
BUF_X1 \mpc/_634_ ( .A(\mpc/_014_ ), .Z(\mpc/_307_ ) );
BUF_X1 \mpc/_635_ ( .A(\mpc/_015_ ), .Z(\mpc/_308_ ) );
BUF_X1 \mpc/_636_ ( .A(\mpc/_016_ ), .Z(\mpc/_309_ ) );
BUF_X1 \mpc/_637_ ( .A(\mpc/_017_ ), .Z(\mpc/_310_ ) );
BUF_X1 \mpc/_638_ ( .A(\mpc/_018_ ), .Z(\mpc/_311_ ) );
BUF_X1 \mpc/_639_ ( .A(\mpc/_019_ ), .Z(\mpc/_312_ ) );
BUF_X1 \mpc/_640_ ( .A(\mpc/_020_ ), .Z(\mpc/_313_ ) );
BUF_X1 \mpc/_641_ ( .A(\mpc/_021_ ), .Z(\mpc/_314_ ) );
BUF_X1 \mpc/_642_ ( .A(\mpc/_022_ ), .Z(\mpc/_315_ ) );
BUF_X1 \mpc/_643_ ( .A(\mpc/_023_ ), .Z(\mpc/_316_ ) );
BUF_X1 \mpc/_644_ ( .A(\mpc/_024_ ), .Z(\mpc/_317_ ) );
BUF_X1 \mpc/_645_ ( .A(\mpc/_025_ ), .Z(\mpc/_318_ ) );
BUF_X1 \mpc/_646_ ( .A(\mpc/_026_ ), .Z(\mpc/_319_ ) );
BUF_X1 \mpc/_647_ ( .A(\mpc/_027_ ), .Z(\mpc/_320_ ) );
BUF_X1 \mpc/_648_ ( .A(\mpc/_028_ ), .Z(\mpc/_321_ ) );
BUF_X1 \mpc/_649_ ( .A(\mpc/_029_ ), .Z(\mpc/_322_ ) );
BUF_X1 \mpc/_650_ ( .A(\mpc/_030_ ), .Z(\mpc/_323_ ) );
BUF_X1 \mpc/_651_ ( .A(\mpc/_031_ ), .Z(\mpc/_324_ ) );
BUF_X1 \mpc/_652_ ( .A(\mpc/_032_ ), .Z(\mpc/_325_ ) );
BUF_X1 \mpc/_653_ ( .A(\mpc/_033_ ), .Z(\mpc/_326_ ) );
INV_X32 \mreg/_06925_ ( .A(\mreg/_03874_ ), .ZN(\mreg/_01055_ ) );
NAND2_X4 \mreg/_06926_ ( .A1(\mreg/_01055_ ), .A2(\mreg/_03873_ ), .ZN(\mreg/_01056_ ) );
INV_X16 \mreg/_06927_ ( .A(\mreg/_03875_ ), .ZN(\mreg/_01057_ ) );
NOR3_X4 \mreg/_06928_ ( .A1(\mreg/_01056_ ), .A2(\mreg/_03876_ ), .A3(\mreg/_01057_ ), .ZN(\mreg/_01058_ ) );
BUF_X4 \mreg/_06929_ ( .A(\mreg/_01058_ ), .Z(\mreg/_01059_ ) );
NAND3_X1 \mreg/_06930_ ( .A1(\mreg/_01059_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04326_ ), .ZN(\mreg/_01060_ ) );
NOR2_X4 \mreg/_06931_ ( .A1(\mreg/_03876_ ), .A2(\mreg/_03875_ ), .ZN(\mreg/_01061_ ) );
BUF_X4 \mreg/_06932_ ( .A(\mreg/_01061_ ), .Z(\mreg/_01062_ ) );
INV_X1 \mreg/_06933_ ( .A(\mreg/_03873_ ), .ZN(\mreg/_01063_ ) );
AND3_X2 \mreg/_06934_ ( .A1(\mreg/_01062_ ), .A2(\mreg/_03874_ ), .A3(\mreg/_01063_ ), .ZN(\mreg/_01064_ ) );
NAND3_X1 \mreg/_06935_ ( .A1(\mreg/_01064_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04198_ ), .ZN(\mreg/_01065_ ) );
AND2_X4 \mreg/_06936_ ( .A1(\mreg/_03874_ ), .A2(\mreg/_03873_ ), .ZN(\mreg/_01066_ ) );
AND2_X4 \mreg/_06937_ ( .A1(\mreg/_01066_ ), .A2(\mreg/_01062_ ), .ZN(\mreg/_01067_ ) );
NAND2_X4 \mreg/_06938_ ( .A1(\mreg/_01067_ ), .A2(\mreg/_03877_ ), .ZN(\mreg/_01068_ ) );
BUF_X4 \mreg/_06939_ ( .A(\mreg/_01068_ ), .Z(\mreg/_01069_ ) );
INV_X1 \mreg/_06940_ ( .A(\mreg/_04230_ ), .ZN(\mreg/_01070_ ) );
OAI21_X1 \mreg/_06941_ ( .A(\mreg/_01065_ ), .B1(\mreg/_01069_ ), .B2(\mreg/_01070_ ), .ZN(\mreg/_01071_ ) );
AND3_X4 \mreg/_06942_ ( .A1(\mreg/_01061_ ), .A2(\mreg/_01055_ ), .A3(\mreg/_03873_ ), .ZN(\mreg/_01072_ ) );
AND2_X1 \mreg/_06943_ ( .A1(\mreg/_01072_ ), .A2(\mreg/_03877_ ), .ZN(\mreg/_01073_ ) );
BUF_X4 \mreg/_06944_ ( .A(\mreg/_01073_ ), .Z(\mreg/_01074_ ) );
BUF_X4 \mreg/_06945_ ( .A(\mreg/_01074_ ), .Z(\mreg/_01075_ ) );
NOR2_X1 \mreg/_06946_ ( .A1(\mreg/_03874_ ), .A2(\mreg/_03873_ ), .ZN(\mreg/_01076_ ) );
AND2_X2 \mreg/_06947_ ( .A1(\mreg/_01076_ ), .A2(\mreg/_03877_ ), .ZN(\mreg/_01077_ ) );
AND2_X1 \mreg/_06948_ ( .A1(\mreg/_01077_ ), .A2(\mreg/_01062_ ), .ZN(\mreg/_01078_ ) );
BUF_X4 \mreg/_06949_ ( .A(\mreg/_01078_ ), .Z(\mreg/_01079_ ) );
BUF_X4 \mreg/_06950_ ( .A(\mreg/_01079_ ), .Z(\mreg/_01080_ ) );
AOI221_X4 \mreg/_06951_ ( .A(\mreg/_01071_ ), .B1(\mreg/_04166_ ), .B2(\mreg/_01075_ ), .C1(\mreg/_04134_ ), .C2(\mreg/_01080_ ), .ZN(\mreg/_01081_ ) );
BUF_X4 \mreg/_06952_ ( .A(\mreg/_01077_ ), .Z(\mreg/_01082_ ) );
BUF_X4 \mreg/_06953_ ( .A(\mreg/_01082_ ), .Z(\mreg/_01083_ ) );
BUF_X4 \mreg/_06954_ ( .A(\mreg/_01083_ ), .Z(\mreg/_01084_ ) );
NOR2_X4 \mreg/_06955_ ( .A1(\mreg/_01057_ ), .A2(\mreg/_03876_ ), .ZN(\mreg/_01085_ ) );
BUF_X4 \mreg/_06956_ ( .A(\mreg/_01085_ ), .Z(\mreg/_01086_ ) );
BUF_X4 \mreg/_06957_ ( .A(\mreg/_01086_ ), .Z(\mreg/_01087_ ) );
NAND3_X1 \mreg/_06958_ ( .A1(\mreg/_01084_ ), .A2(\mreg/_04294_ ), .A3(\mreg/_01087_ ), .ZN(\mreg/_01088_ ) );
NOR2_X4 \mreg/_06959_ ( .A1(\mreg/_01055_ ), .A2(\mreg/_03873_ ), .ZN(\mreg/_01089_ ) );
AND2_X4 \mreg/_06960_ ( .A1(\mreg/_01089_ ), .A2(\mreg/_01085_ ), .ZN(\mreg/_01090_ ) );
BUF_X4 \mreg/_06961_ ( .A(\mreg/_01090_ ), .Z(\mreg/_01091_ ) );
BUF_X4 \mreg/_06962_ ( .A(\mreg/_01091_ ), .Z(\mreg/_01092_ ) );
NAND3_X1 \mreg/_06963_ ( .A1(\mreg/_01092_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04358_ ), .ZN(\mreg/_01093_ ) );
INV_X32 \mreg/_06964_ ( .A(\mreg/_03876_ ), .ZN(\mreg/_01094_ ) );
AND3_X4 \mreg/_06965_ ( .A1(\mreg/_01066_ ), .A2(\mreg/_01094_ ), .A3(\mreg/_03875_ ), .ZN(\mreg/_01095_ ) );
BUF_X8 \mreg/_06966_ ( .A(\mreg/_01095_ ), .Z(\mreg/_01096_ ) );
BUF_X8 \mreg/_06967_ ( .A(\mreg/_01096_ ), .Z(\mreg/_01097_ ) );
BUF_X2 \mreg/_06968_ ( .A(\mreg/_01097_ ), .Z(\mreg/_01098_ ) );
NAND3_X1 \mreg/_06969_ ( .A1(\mreg/_01098_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04390_ ), .ZN(\mreg/_01099_ ) );
AND2_X1 \mreg/_06970_ ( .A1(\mreg/_01093_ ), .A2(\mreg/_01099_ ), .ZN(\mreg/_01100_ ) );
AND4_X1 \mreg/_06971_ ( .A1(\mreg/_01060_ ), .A2(\mreg/_01081_ ), .A3(\mreg/_01088_ ), .A4(\mreg/_01100_ ), .ZN(\mreg/_01101_ ) );
INV_X1 \mreg/_06972_ ( .A(\mreg/_03877_ ), .ZN(\mreg/_01102_ ) );
CLKBUF_X2 \mreg/_06973_ ( .A(\mreg/_01102_ ), .Z(\mreg/_01103_ ) );
AND3_X1 \mreg/_06974_ ( .A1(\mreg/_01064_ ), .A2(\mreg/_01103_ ), .A3(\mreg/_04614_ ), .ZN(\mreg/_01104_ ) );
AND2_X4 \mreg/_06975_ ( .A1(\mreg/_01067_ ), .A2(\mreg/_01102_ ), .ZN(\mreg/_01105_ ) );
BUF_X4 \mreg/_06976_ ( .A(\mreg/_01105_ ), .Z(\mreg/_01106_ ) );
BUF_X2 \mreg/_06977_ ( .A(\mreg/_01072_ ), .Z(\mreg/_01107_ ) );
BUF_X4 \mreg/_06978_ ( .A(\mreg/_01102_ ), .Z(\mreg/_01108_ ) );
BUF_X2 \mreg/_06979_ ( .A(\mreg/_01108_ ), .Z(\mreg/_01109_ ) );
AND2_X1 \mreg/_06980_ ( .A1(\mreg/_01107_ ), .A2(\mreg/_01109_ ), .ZN(\mreg/_01110_ ) );
AOI221_X4 \mreg/_06981_ ( .A(\mreg/_01104_ ), .B1(\mreg/_01106_ ), .B2(\mreg/_04710_ ), .C1(\mreg/_04262_ ), .C2(\mreg/_01110_ ), .ZN(\mreg/_01111_ ) );
AND3_X2 \mreg/_06982_ ( .A1(\mreg/_01066_ ), .A2(\mreg/_03876_ ), .A3(\mreg/_01057_ ), .ZN(\mreg/_01112_ ) );
BUF_X4 \mreg/_06983_ ( .A(\mreg/_01112_ ), .Z(\mreg/_01113_ ) );
BUF_X2 \mreg/_06984_ ( .A(\mreg/_01109_ ), .Z(\mreg/_01114_ ) );
AND3_X1 \mreg/_06985_ ( .A1(\mreg/_01113_ ), .A2(\mreg/_01114_ ), .A3(\mreg/_03974_ ), .ZN(\mreg/_01115_ ) );
NOR2_X2 \mreg/_06986_ ( .A1(\mreg/_01094_ ), .A2(\mreg/_03875_ ), .ZN(\mreg/_01116_ ) );
AND2_X4 \mreg/_06987_ ( .A1(\mreg/_01089_ ), .A2(\mreg/_01116_ ), .ZN(\mreg/_01117_ ) );
BUF_X2 \mreg/_06988_ ( .A(\mreg/_01103_ ), .Z(\mreg/_01118_ ) );
AND3_X1 \mreg/_06989_ ( .A1(\mreg/_01117_ ), .A2(\mreg/_01118_ ), .A3(\mreg/_03942_ ), .ZN(\mreg/_01119_ ) );
NOR3_X1 \mreg/_06990_ ( .A1(\mreg/_01056_ ), .A2(\mreg/_01094_ ), .A3(\mreg/_03875_ ), .ZN(\mreg/_01120_ ) );
BUF_X2 \mreg/_06991_ ( .A(\mreg/_01120_ ), .Z(\mreg/_01121_ ) );
BUF_X2 \mreg/_06992_ ( .A(\mreg/_01108_ ), .Z(\mreg/_01122_ ) );
AND3_X1 \mreg/_06993_ ( .A1(\mreg/_01121_ ), .A2(\mreg/_01122_ ), .A3(\mreg/_04902_ ), .ZN(\mreg/_01123_ ) );
NOR3_X1 \mreg/_06994_ ( .A1(\mreg/_03877_ ), .A2(\mreg/_03874_ ), .A3(\mreg/_03873_ ), .ZN(\mreg/_01124_ ) );
BUF_X4 \mreg/_06995_ ( .A(\mreg/_01124_ ), .Z(\mreg/_01125_ ) );
BUF_X2 \mreg/_06996_ ( .A(\mreg/_01125_ ), .Z(\mreg/_01126_ ) );
CLKBUF_X2 \mreg/_06997_ ( .A(\mreg/_01116_ ), .Z(\mreg/_01127_ ) );
AND3_X1 \mreg/_06998_ ( .A1(\mreg/_01126_ ), .A2(\mreg/_04870_ ), .A3(\mreg/_01127_ ), .ZN(\mreg/_01128_ ) );
NOR4_X1 \mreg/_06999_ ( .A1(\mreg/_01115_ ), .A2(\mreg/_01119_ ), .A3(\mreg/_01123_ ), .A4(\mreg/_01128_ ), .ZN(\mreg/_01129_ ) );
BUF_X4 \mreg/_07000_ ( .A(\mreg/_01122_ ), .Z(\mreg/_01130_ ) );
NAND3_X1 \mreg/_07001_ ( .A1(\mreg/_01092_ ), .A2(\mreg/_01130_ ), .A3(\mreg/_04806_ ), .ZN(\mreg/_01131_ ) );
NAND3_X1 \mreg/_07002_ ( .A1(\mreg/_01098_ ), .A2(\mreg/_01114_ ), .A3(\mreg/_04838_ ), .ZN(\mreg/_01132_ ) );
CLKBUF_X2 \mreg/_07003_ ( .A(\mreg/_01109_ ), .Z(\mreg/_01133_ ) );
NAND3_X1 \mreg/_07004_ ( .A1(\mreg/_01058_ ), .A2(\mreg/_01133_ ), .A3(\mreg/_04774_ ), .ZN(\mreg/_01134_ ) );
NAND3_X1 \mreg/_07005_ ( .A1(\mreg/_01126_ ), .A2(\mreg/_01086_ ), .A3(\mreg/_04742_ ), .ZN(\mreg/_01135_ ) );
AND4_X1 \mreg/_07006_ ( .A1(\mreg/_01131_ ), .A2(\mreg/_01132_ ), .A3(\mreg/_01134_ ), .A4(\mreg/_01135_ ), .ZN(\mreg/_01136_ ) );
AND2_X4 \mreg/_07007_ ( .A1(\mreg/_03876_ ), .A2(\mreg/_03875_ ), .ZN(\mreg/_01137_ ) );
AND2_X4 \mreg/_07008_ ( .A1(\mreg/_01066_ ), .A2(\mreg/_01137_ ), .ZN(\mreg/_01138_ ) );
BUF_X8 \mreg/_07009_ ( .A(\mreg/_01138_ ), .Z(\mreg/_01139_ ) );
BUF_X4 \mreg/_07010_ ( .A(\mreg/_01139_ ), .Z(\mreg/_01140_ ) );
NAND3_X1 \mreg/_07011_ ( .A1(\mreg/_01140_ ), .A2(\mreg/_01130_ ), .A3(\mreg/_04102_ ), .ZN(\mreg/_01141_ ) );
AND3_X2 \mreg/_07012_ ( .A1(\mreg/_01137_ ), .A2(\mreg/_03874_ ), .A3(\mreg/_01063_ ), .ZN(\mreg/_01142_ ) );
BUF_X2 \mreg/_07013_ ( .A(\mreg/_01142_ ), .Z(\mreg/_01143_ ) );
BUF_X2 \mreg/_07014_ ( .A(\mreg/_01109_ ), .Z(\mreg/_01144_ ) );
NAND3_X1 \mreg/_07015_ ( .A1(\mreg/_01143_ ), .A2(\mreg/_01144_ ), .A3(\mreg/_04070_ ), .ZN(\mreg/_01145_ ) );
NOR3_X1 \mreg/_07016_ ( .A1(\mreg/_01056_ ), .A2(\mreg/_01094_ ), .A3(\mreg/_01057_ ), .ZN(\mreg/_01146_ ) );
BUF_X4 \mreg/_07017_ ( .A(\mreg/_01146_ ), .Z(\mreg/_01147_ ) );
BUF_X2 \mreg/_07018_ ( .A(\mreg/_01147_ ), .Z(\mreg/_01148_ ) );
NAND3_X1 \mreg/_07019_ ( .A1(\mreg/_01148_ ), .A2(\mreg/_01133_ ), .A3(\mreg/_04038_ ), .ZN(\mreg/_01149_ ) );
BUF_X4 \mreg/_07020_ ( .A(\mreg/_01137_ ), .Z(\mreg/_01150_ ) );
BUF_X2 \mreg/_07021_ ( .A(\mreg/_01150_ ), .Z(\mreg/_01151_ ) );
NAND3_X1 \mreg/_07022_ ( .A1(\mreg/_01126_ ), .A2(\mreg/_04006_ ), .A3(\mreg/_01151_ ), .ZN(\mreg/_01152_ ) );
AND4_X1 \mreg/_07023_ ( .A1(\mreg/_01141_ ), .A2(\mreg/_01145_ ), .A3(\mreg/_01149_ ), .A4(\mreg/_01152_ ), .ZN(\mreg/_01153_ ) );
AND4_X1 \mreg/_07024_ ( .A1(\mreg/_01111_ ), .A2(\mreg/_01129_ ), .A3(\mreg/_01136_ ), .A4(\mreg/_01153_ ), .ZN(\mreg/_01154_ ) );
BUF_X2 \mreg/_07025_ ( .A(\mreg/_01121_ ), .Z(\mreg/_01155_ ) );
BUF_X4 \mreg/_07026_ ( .A(\mreg/_01155_ ), .Z(\mreg/_01156_ ) );
NAND3_X1 \mreg/_07027_ ( .A1(\mreg/_01156_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04454_ ), .ZN(\mreg/_01157_ ) );
BUF_X4 \mreg/_07028_ ( .A(\mreg/_01117_ ), .Z(\mreg/_01158_ ) );
BUF_X4 \mreg/_07029_ ( .A(\mreg/_01158_ ), .Z(\mreg/_01159_ ) );
NAND3_X1 \mreg/_07030_ ( .A1(\mreg/_01159_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04486_ ), .ZN(\mreg/_01160_ ) );
BUF_X4 \mreg/_07031_ ( .A(\mreg/_01116_ ), .Z(\mreg/_01161_ ) );
BUF_X2 \mreg/_07032_ ( .A(\mreg/_01161_ ), .Z(\mreg/_01162_ ) );
BUF_X2 \mreg/_07033_ ( .A(\mreg/_01162_ ), .Z(\mreg/_01163_ ) );
NAND3_X1 \mreg/_07034_ ( .A1(\mreg/_01084_ ), .A2(\mreg/_04422_ ), .A3(\mreg/_01163_ ), .ZN(\mreg/_01164_ ) );
BUF_X4 \mreg/_07035_ ( .A(\mreg/_01113_ ), .Z(\mreg/_01165_ ) );
NAND3_X1 \mreg/_07036_ ( .A1(\mreg/_01165_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04518_ ), .ZN(\mreg/_01166_ ) );
AND4_X1 \mreg/_07037_ ( .A1(\mreg/_01157_ ), .A2(\mreg/_01160_ ), .A3(\mreg/_01164_ ), .A4(\mreg/_01166_ ), .ZN(\mreg/_01167_ ) );
NAND3_X1 \mreg/_07038_ ( .A1(\mreg/_01147_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04582_ ), .ZN(\mreg/_01168_ ) );
NAND3_X1 \mreg/_07039_ ( .A1(\mreg/_01082_ ), .A2(\mreg/_04550_ ), .A3(\mreg/_01151_ ), .ZN(\mreg/_01169_ ) );
NAND2_X1 \mreg/_07040_ ( .A1(\mreg/_01168_ ), .A2(\mreg/_01169_ ), .ZN(\mreg/_01170_ ) );
AND2_X4 \mreg/_07041_ ( .A1(\mreg/_01139_ ), .A2(\mreg/_03877_ ), .ZN(\mreg/_01171_ ) );
BUF_X8 \mreg/_07042_ ( .A(\mreg/_01171_ ), .Z(\mreg/_01172_ ) );
BUF_X4 \mreg/_07043_ ( .A(\mreg/_01172_ ), .Z(\mreg/_01173_ ) );
AND2_X2 \mreg/_07044_ ( .A1(\mreg/_01142_ ), .A2(\mreg/_03877_ ), .ZN(\mreg/_01174_ ) );
BUF_X4 \mreg/_07045_ ( .A(\mreg/_01174_ ), .Z(\mreg/_01175_ ) );
AOI221_X4 \mreg/_07046_ ( .A(\mreg/_01170_ ), .B1(\mreg/_04678_ ), .B2(\mreg/_01173_ ), .C1(\mreg/_04646_ ), .C2(\mreg/_01175_ ), .ZN(\mreg/_01176_ ) );
NAND4_X1 \mreg/_07047_ ( .A1(\mreg/_01101_ ), .A2(\mreg/_01154_ ), .A3(\mreg/_01167_ ), .A4(\mreg/_01176_ ), .ZN(\mreg/_03910_ ) );
BUF_X4 \mreg/_07048_ ( .A(\mreg/_01082_ ), .Z(\mreg/_01177_ ) );
BUF_X4 \mreg/_07049_ ( .A(\mreg/_01150_ ), .Z(\mreg/_01178_ ) );
NAND3_X1 \mreg/_07050_ ( .A1(\mreg/_01177_ ), .A2(\mreg/_04561_ ), .A3(\mreg/_01178_ ), .ZN(\mreg/_01179_ ) );
BUF_X4 \mreg/_07051_ ( .A(\mreg/_01142_ ), .Z(\mreg/_01180_ ) );
NAND3_X1 \mreg/_07052_ ( .A1(\mreg/_01180_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04657_ ), .ZN(\mreg/_01181_ ) );
BUF_X4 \mreg/_07053_ ( .A(\mreg/_01147_ ), .Z(\mreg/_01182_ ) );
NAND3_X1 \mreg/_07054_ ( .A1(\mreg/_01182_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04593_ ), .ZN(\mreg/_01183_ ) );
BUF_X4 \mreg/_07055_ ( .A(\mreg/_01139_ ), .Z(\mreg/_01184_ ) );
INV_X1 \mreg/_07056_ ( .A(\mreg/_00031_ ), .ZN(\mreg/_01185_ ) );
NAND3_X1 \mreg/_07057_ ( .A1(\mreg/_01184_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_01185_ ), .ZN(\mreg/_01186_ ) );
AND4_X1 \mreg/_07058_ ( .A1(\mreg/_01179_ ), .A2(\mreg/_01181_ ), .A3(\mreg/_01183_ ), .A4(\mreg/_01186_ ), .ZN(\mreg/_01187_ ) );
BUF_X4 \mreg/_07059_ ( .A(\mreg/_01089_ ), .Z(\mreg/_01188_ ) );
NAND4_X1 \mreg/_07060_ ( .A1(\mreg/_01188_ ), .A2(\mreg/_01161_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04497_ ), .ZN(\mreg/_01189_ ) );
NAND2_X4 \mreg/_07061_ ( .A1(\mreg/_01112_ ), .A2(\mreg/_03877_ ), .ZN(\mreg/_01190_ ) );
BUF_X4 \mreg/_07062_ ( .A(\mreg/_01190_ ), .Z(\mreg/_01191_ ) );
INV_X1 \mreg/_07063_ ( .A(\mreg/_04529_ ), .ZN(\mreg/_01192_ ) );
OAI21_X1 \mreg/_07064_ ( .A(\mreg/_01189_ ), .B1(\mreg/_01191_ ), .B2(\mreg/_01192_ ), .ZN(\mreg/_01193_ ) );
AND2_X1 \mreg/_07065_ ( .A1(\mreg/_01120_ ), .A2(\mreg/_03877_ ), .ZN(\mreg/_01194_ ) );
BUF_X4 \mreg/_07066_ ( .A(\mreg/_01194_ ), .Z(\mreg/_01195_ ) );
BUF_X4 \mreg/_07067_ ( .A(\mreg/_01195_ ), .Z(\mreg/_01196_ ) );
AND2_X1 \mreg/_07068_ ( .A1(\mreg/_01077_ ), .A2(\mreg/_01116_ ), .ZN(\mreg/_01197_ ) );
BUF_X4 \mreg/_07069_ ( .A(\mreg/_01197_ ), .Z(\mreg/_01198_ ) );
AOI221_X4 \mreg/_07070_ ( .A(\mreg/_01193_ ), .B1(\mreg/_04465_ ), .B2(\mreg/_01196_ ), .C1(\mreg/_04433_ ), .C2(\mreg/_01198_ ), .ZN(\mreg/_01199_ ) );
NAND3_X1 \mreg/_07071_ ( .A1(\mreg/_01091_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04369_ ), .ZN(\mreg/_01200_ ) );
NAND3_X1 \mreg/_07072_ ( .A1(\mreg/_01097_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04401_ ), .ZN(\mreg/_01201_ ) );
NAND2_X1 \mreg/_07073_ ( .A1(\mreg/_01200_ ), .A2(\mreg/_01201_ ), .ZN(\mreg/_01202_ ) );
AND2_X4 \mreg/_07074_ ( .A1(\mreg/_01058_ ), .A2(\mreg/_03877_ ), .ZN(\mreg/_01203_ ) );
BUF_X4 \mreg/_07075_ ( .A(\mreg/_01203_ ), .Z(\mreg/_01204_ ) );
BUF_X4 \mreg/_07076_ ( .A(\mreg/_01204_ ), .Z(\mreg/_01205_ ) );
AND2_X2 \mreg/_07077_ ( .A1(\mreg/_01077_ ), .A2(\mreg/_01085_ ), .ZN(\mreg/_01206_ ) );
BUF_X4 \mreg/_07078_ ( .A(\mreg/_01206_ ), .Z(\mreg/_01207_ ) );
AOI221_X4 \mreg/_07079_ ( .A(\mreg/_01202_ ), .B1(\mreg/_04337_ ), .B2(\mreg/_01205_ ), .C1(\mreg/_04305_ ), .C2(\mreg/_01207_ ), .ZN(\mreg/_01208_ ) );
BUF_X4 \mreg/_07080_ ( .A(\mreg/_01062_ ), .Z(\mreg/_01209_ ) );
NAND4_X1 \mreg/_07081_ ( .A1(\mreg/_01188_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04209_ ), .A4(\mreg/_01209_ ), .ZN(\mreg/_01210_ ) );
BUF_X4 \mreg/_07082_ ( .A(\mreg/_01066_ ), .Z(\mreg/_01211_ ) );
BUF_X4 \mreg/_07083_ ( .A(\mreg/_01062_ ), .Z(\mreg/_01212_ ) );
NAND4_X1 \mreg/_07084_ ( .A1(\mreg/_01211_ ), .A2(\mreg/_01212_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04241_ ), .ZN(\mreg/_01213_ ) );
NAND2_X1 \mreg/_07085_ ( .A1(\mreg/_01210_ ), .A2(\mreg/_01213_ ), .ZN(\mreg/_01214_ ) );
AOI221_X4 \mreg/_07086_ ( .A(\mreg/_01214_ ), .B1(\mreg/_04177_ ), .B2(\mreg/_01075_ ), .C1(\mreg/_04145_ ), .C2(\mreg/_01080_ ), .ZN(\mreg/_01215_ ) );
AND4_X2 \mreg/_07087_ ( .A1(\mreg/_01187_ ), .A2(\mreg/_01199_ ), .A3(\mreg/_01208_ ), .A4(\mreg/_01215_ ), .ZN(\mreg/_01216_ ) );
BUF_X2 \mreg/_07088_ ( .A(\mreg/_01109_ ), .Z(\mreg/_01217_ ) );
AND3_X1 \mreg/_07089_ ( .A1(\mreg/_01107_ ), .A2(\mreg/_01217_ ), .A3(\mreg/_04273_ ), .ZN(\mreg/_01218_ ) );
BUF_X4 \mreg/_07090_ ( .A(\mreg/_01105_ ), .Z(\mreg/_01219_ ) );
AND2_X1 \mreg/_07091_ ( .A1(\mreg/_01064_ ), .A2(\mreg/_01102_ ), .ZN(\mreg/_01220_ ) );
BUF_X4 \mreg/_07092_ ( .A(\mreg/_01220_ ), .Z(\mreg/_01221_ ) );
BUF_X4 \mreg/_07093_ ( .A(\mreg/_01221_ ), .Z(\mreg/_01222_ ) );
AOI221_X4 \mreg/_07094_ ( .A(\mreg/_01218_ ), .B1(\mreg/_01219_ ), .B2(\mreg/_04721_ ), .C1(\mreg/_04625_ ), .C2(\mreg/_01222_ ), .ZN(\mreg/_01223_ ) );
AND3_X1 \mreg/_07095_ ( .A1(\mreg/_01091_ ), .A2(\mreg/_01109_ ), .A3(\mreg/_04817_ ), .ZN(\mreg/_01224_ ) );
AND3_X1 \mreg/_07096_ ( .A1(\mreg/_01097_ ), .A2(\mreg/_01109_ ), .A3(\mreg/_04849_ ), .ZN(\mreg/_01225_ ) );
OR2_X1 \mreg/_07097_ ( .A1(\mreg/_01224_ ), .A2(\mreg/_01225_ ), .ZN(\mreg/_01226_ ) );
AND2_X1 \mreg/_07098_ ( .A1(\mreg/_01058_ ), .A2(\mreg/_01108_ ), .ZN(\mreg/_01227_ ) );
BUF_X4 \mreg/_07099_ ( .A(\mreg/_01227_ ), .Z(\mreg/_01228_ ) );
AND2_X2 \mreg/_07100_ ( .A1(\mreg/_01124_ ), .A2(\mreg/_01085_ ), .ZN(\mreg/_01229_ ) );
BUF_X4 \mreg/_07101_ ( .A(\mreg/_01229_ ), .Z(\mreg/_01230_ ) );
AOI221_X4 \mreg/_07102_ ( .A(\mreg/_01226_ ), .B1(\mreg/_04785_ ), .B2(\mreg/_01228_ ), .C1(\mreg/_04753_ ), .C2(\mreg/_01230_ ), .ZN(\mreg/_01231_ ) );
BUF_X2 \mreg/_07103_ ( .A(\mreg/_01142_ ), .Z(\mreg/_01232_ ) );
CLKBUF_X2 \mreg/_07104_ ( .A(\mreg/_01118_ ), .Z(\mreg/_01233_ ) );
NAND3_X1 \mreg/_07105_ ( .A1(\mreg/_01232_ ), .A2(\mreg/_01233_ ), .A3(\mreg/_04081_ ), .ZN(\mreg/_01234_ ) );
BUF_X2 \mreg/_07106_ ( .A(\mreg/_01147_ ), .Z(\mreg/_01235_ ) );
BUF_X2 \mreg/_07107_ ( .A(\mreg/_01118_ ), .Z(\mreg/_01236_ ) );
NAND3_X1 \mreg/_07108_ ( .A1(\mreg/_01235_ ), .A2(\mreg/_01236_ ), .A3(\mreg/_04049_ ), .ZN(\mreg/_01237_ ) );
BUF_X2 \mreg/_07109_ ( .A(\mreg/_01140_ ), .Z(\mreg/_01238_ ) );
BUF_X2 \mreg/_07110_ ( .A(\mreg/_01118_ ), .Z(\mreg/_01239_ ) );
NAND3_X1 \mreg/_07111_ ( .A1(\mreg/_01238_ ), .A2(\mreg/_01239_ ), .A3(\mreg/_04113_ ), .ZN(\mreg/_01240_ ) );
BUF_X2 \mreg/_07112_ ( .A(\mreg/_01126_ ), .Z(\mreg/_01241_ ) );
BUF_X2 \mreg/_07113_ ( .A(\mreg/_01151_ ), .Z(\mreg/_01242_ ) );
NAND3_X1 \mreg/_07114_ ( .A1(\mreg/_01241_ ), .A2(\mreg/_04017_ ), .A3(\mreg/_01242_ ), .ZN(\mreg/_01243_ ) );
NAND4_X1 \mreg/_07115_ ( .A1(\mreg/_01234_ ), .A2(\mreg/_01237_ ), .A3(\mreg/_01240_ ), .A4(\mreg/_01243_ ), .ZN(\mreg/_01244_ ) );
NAND3_X1 \mreg/_07116_ ( .A1(\mreg/_01158_ ), .A2(\mreg/_01236_ ), .A3(\mreg/_03953_ ), .ZN(\mreg/_01245_ ) );
NAND3_X1 \mreg/_07117_ ( .A1(\mreg/_01113_ ), .A2(\mreg/_01236_ ), .A3(\mreg/_03985_ ), .ZN(\mreg/_01246_ ) );
NAND2_X1 \mreg/_07118_ ( .A1(\mreg/_01245_ ), .A2(\mreg/_01246_ ), .ZN(\mreg/_01247_ ) );
CLKBUF_X2 \mreg/_07119_ ( .A(\mreg/_01122_ ), .Z(\mreg/_01248_ ) );
AND3_X1 \mreg/_07120_ ( .A1(\mreg/_01155_ ), .A2(\mreg/_01248_ ), .A3(\mreg/_04913_ ), .ZN(\mreg/_01249_ ) );
CLKBUF_X2 \mreg/_07121_ ( .A(\mreg/_01126_ ), .Z(\mreg/_01250_ ) );
BUF_X2 \mreg/_07122_ ( .A(\mreg/_01127_ ), .Z(\mreg/_01251_ ) );
AND3_X1 \mreg/_07123_ ( .A1(\mreg/_01250_ ), .A2(\mreg/_04881_ ), .A3(\mreg/_01251_ ), .ZN(\mreg/_01252_ ) );
NOR4_X1 \mreg/_07124_ ( .A1(\mreg/_01244_ ), .A2(\mreg/_01247_ ), .A3(\mreg/_01249_ ), .A4(\mreg/_01252_ ), .ZN(\mreg/_01253_ ) );
NAND4_X1 \mreg/_07125_ ( .A1(\mreg/_01216_ ), .A2(\mreg/_01223_ ), .A3(\mreg/_01231_ ), .A4(\mreg/_01253_ ), .ZN(\mreg/_03921_ ) );
NAND3_X1 \mreg/_07126_ ( .A1(\mreg/_01147_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04604_ ), .ZN(\mreg/_01254_ ) );
BUF_X2 \mreg/_07127_ ( .A(\mreg/_01077_ ), .Z(\mreg/_01255_ ) );
NAND3_X1 \mreg/_07128_ ( .A1(\mreg/_01255_ ), .A2(\mreg/_04572_ ), .A3(\mreg/_01150_ ), .ZN(\mreg/_01256_ ) );
NAND2_X1 \mreg/_07129_ ( .A1(\mreg/_01254_ ), .A2(\mreg/_01256_ ), .ZN(\mreg/_01257_ ) );
INV_X1 \mreg/_07130_ ( .A(\mreg/_00032_ ), .ZN(\mreg/_01258_ ) );
AOI221_X1 \mreg/_07131_ ( .A(\mreg/_01257_ ), .B1(\mreg/_01258_ ), .B2(\mreg/_01173_ ), .C1(\mreg/_04668_ ), .C2(\mreg/_01175_ ), .ZN(\mreg/_01259_ ) );
AND3_X1 \mreg/_07132_ ( .A1(\mreg/_01077_ ), .A2(\mreg/_04444_ ), .A3(\mreg/_01127_ ), .ZN(\mreg/_01260_ ) );
NAND4_X1 \mreg/_07133_ ( .A1(\mreg/_01188_ ), .A2(\mreg/_01161_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04508_ ), .ZN(\mreg/_01261_ ) );
INV_X1 \mreg/_07134_ ( .A(\mreg/_04540_ ), .ZN(\mreg/_01262_ ) );
OAI21_X1 \mreg/_07135_ ( .A(\mreg/_01261_ ), .B1(\mreg/_01191_ ), .B2(\mreg/_01262_ ), .ZN(\mreg/_01263_ ) );
AOI211_X4 \mreg/_07136_ ( .A(\mreg/_01260_ ), .B(\mreg/_01263_ ), .C1(\mreg/_04476_ ), .C2(\mreg/_01196_ ), .ZN(\mreg/_01264_ ) );
NAND3_X1 \mreg/_07137_ ( .A1(\mreg/_01091_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04380_ ), .ZN(\mreg/_01265_ ) );
NAND3_X1 \mreg/_07138_ ( .A1(\mreg/_01097_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04412_ ), .ZN(\mreg/_01266_ ) );
NAND2_X1 \mreg/_07139_ ( .A1(\mreg/_01265_ ), .A2(\mreg/_01266_ ), .ZN(\mreg/_01267_ ) );
AOI221_X4 \mreg/_07140_ ( .A(\mreg/_01267_ ), .B1(\mreg/_04348_ ), .B2(\mreg/_01205_ ), .C1(\mreg/_04316_ ), .C2(\mreg/_01207_ ), .ZN(\mreg/_01268_ ) );
BUF_X4 \mreg/_07141_ ( .A(\mreg/_01089_ ), .Z(\mreg/_01269_ ) );
NAND4_X1 \mreg/_07142_ ( .A1(\mreg/_01269_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04220_ ), .A4(\mreg/_01209_ ), .ZN(\mreg/_01270_ ) );
INV_X1 \mreg/_07143_ ( .A(\mreg/_04252_ ), .ZN(\mreg/_01271_ ) );
OAI21_X1 \mreg/_07144_ ( .A(\mreg/_01270_ ), .B1(\mreg/_01069_ ), .B2(\mreg/_01271_ ), .ZN(\mreg/_01272_ ) );
AOI221_X4 \mreg/_07145_ ( .A(\mreg/_01272_ ), .B1(\mreg/_04188_ ), .B2(\mreg/_01075_ ), .C1(\mreg/_04156_ ), .C2(\mreg/_01080_ ), .ZN(\mreg/_01273_ ) );
AND4_X4 \mreg/_07146_ ( .A1(\mreg/_01259_ ), .A2(\mreg/_01264_ ), .A3(\mreg/_01268_ ), .A4(\mreg/_01273_ ), .ZN(\mreg/_01274_ ) );
BUF_X4 \mreg/_07147_ ( .A(\mreg/_01092_ ), .Z(\mreg/_01275_ ) );
BUF_X4 \mreg/_07148_ ( .A(\mreg/_01122_ ), .Z(\mreg/_01276_ ) );
BUF_X4 \mreg/_07149_ ( .A(\mreg/_01276_ ), .Z(\mreg/_01277_ ) );
NAND3_X1 \mreg/_07150_ ( .A1(\mreg/_01275_ ), .A2(\mreg/_01277_ ), .A3(\mreg/_04828_ ), .ZN(\mreg/_01278_ ) );
AND3_X1 \mreg/_07151_ ( .A1(\mreg/_01072_ ), .A2(\mreg/_01103_ ), .A3(\mreg/_04284_ ), .ZN(\mreg/_01279_ ) );
AOI221_X4 \mreg/_07152_ ( .A(\mreg/_01279_ ), .B1(\mreg/_01106_ ), .B2(\mreg/_04732_ ), .C1(\mreg/_04636_ ), .C2(\mreg/_01221_ ), .ZN(\mreg/_01280_ ) );
BUF_X4 \mreg/_07153_ ( .A(\mreg/_01098_ ), .Z(\mreg/_01281_ ) );
BUF_X4 \mreg/_07154_ ( .A(\mreg/_01276_ ), .Z(\mreg/_01282_ ) );
NAND3_X1 \mreg/_07155_ ( .A1(\mreg/_01281_ ), .A2(\mreg/_01282_ ), .A3(\mreg/_04860_ ), .ZN(\mreg/_01283_ ) );
BUF_X4 \mreg/_07156_ ( .A(\mreg/_01228_ ), .Z(\mreg/_01284_ ) );
AOI22_X1 \mreg/_07157_ ( .A1(\mreg/_01284_ ), .A2(\mreg/_04796_ ), .B1(\mreg/_04764_ ), .B2(\mreg/_01230_ ), .ZN(\mreg/_01285_ ) );
AND4_X1 \mreg/_07158_ ( .A1(\mreg/_01278_ ), .A2(\mreg/_01280_ ), .A3(\mreg/_01283_ ), .A4(\mreg/_01285_ ), .ZN(\mreg/_01286_ ) );
BUF_X4 \mreg/_07159_ ( .A(\mreg/_01276_ ), .Z(\mreg/_01287_ ) );
NAND3_X1 \mreg/_07160_ ( .A1(\mreg/_01156_ ), .A2(\mreg/_01287_ ), .A3(\mreg/_04924_ ), .ZN(\mreg/_01288_ ) );
BUF_X4 \mreg/_07161_ ( .A(\mreg/_01276_ ), .Z(\mreg/_01289_ ) );
NAND3_X1 \mreg/_07162_ ( .A1(\mreg/_01159_ ), .A2(\mreg/_01289_ ), .A3(\mreg/_03964_ ), .ZN(\mreg/_01290_ ) );
BUF_X4 \mreg/_07163_ ( .A(\mreg/_01125_ ), .Z(\mreg/_01291_ ) );
BUF_X4 \mreg/_07164_ ( .A(\mreg/_01291_ ), .Z(\mreg/_01292_ ) );
BUF_X4 \mreg/_07165_ ( .A(\mreg/_01251_ ), .Z(\mreg/_01293_ ) );
NAND3_X1 \mreg/_07166_ ( .A1(\mreg/_01292_ ), .A2(\mreg/_01293_ ), .A3(\mreg/_04892_ ), .ZN(\mreg/_01294_ ) );
BUF_X4 \mreg/_07167_ ( .A(\mreg/_01276_ ), .Z(\mreg/_01295_ ) );
NAND3_X1 \mreg/_07168_ ( .A1(\mreg/_01165_ ), .A2(\mreg/_01295_ ), .A3(\mreg/_03996_ ), .ZN(\mreg/_01296_ ) );
AND4_X1 \mreg/_07169_ ( .A1(\mreg/_01288_ ), .A2(\mreg/_01290_ ), .A3(\mreg/_01294_ ), .A4(\mreg/_01296_ ), .ZN(\mreg/_01297_ ) );
BUF_X4 \mreg/_07170_ ( .A(\mreg/_01291_ ), .Z(\mreg/_01298_ ) );
BUF_X4 \mreg/_07171_ ( .A(\mreg/_01178_ ), .Z(\mreg/_01299_ ) );
NAND3_X1 \mreg/_07172_ ( .A1(\mreg/_01298_ ), .A2(\mreg/_04028_ ), .A3(\mreg/_01299_ ), .ZN(\mreg/_01300_ ) );
BUF_X4 \mreg/_07173_ ( .A(\mreg/_01180_ ), .Z(\mreg/_01301_ ) );
BUF_X4 \mreg/_07174_ ( .A(\mreg/_01276_ ), .Z(\mreg/_01302_ ) );
NAND3_X1 \mreg/_07175_ ( .A1(\mreg/_01301_ ), .A2(\mreg/_01302_ ), .A3(\mreg/_04092_ ), .ZN(\mreg/_01303_ ) );
BUF_X4 \mreg/_07176_ ( .A(\mreg/_01147_ ), .Z(\mreg/_01304_ ) );
BUF_X4 \mreg/_07177_ ( .A(\mreg/_01304_ ), .Z(\mreg/_01305_ ) );
BUF_X4 \mreg/_07178_ ( .A(\mreg/_01276_ ), .Z(\mreg/_01306_ ) );
NAND3_X1 \mreg/_07179_ ( .A1(\mreg/_01305_ ), .A2(\mreg/_01306_ ), .A3(\mreg/_04060_ ), .ZN(\mreg/_01307_ ) );
BUF_X4 \mreg/_07180_ ( .A(\mreg/_01184_ ), .Z(\mreg/_01308_ ) );
BUF_X2 \mreg/_07181_ ( .A(\mreg/_01130_ ), .Z(\mreg/_01309_ ) );
NAND3_X1 \mreg/_07182_ ( .A1(\mreg/_01308_ ), .A2(\mreg/_01309_ ), .A3(\mreg/_04124_ ), .ZN(\mreg/_01310_ ) );
AND4_X1 \mreg/_07183_ ( .A1(\mreg/_01300_ ), .A2(\mreg/_01303_ ), .A3(\mreg/_01307_ ), .A4(\mreg/_01310_ ), .ZN(\mreg/_01311_ ) );
NAND4_X1 \mreg/_07184_ ( .A1(\mreg/_01274_ ), .A2(\mreg/_01286_ ), .A3(\mreg/_01297_ ), .A4(\mreg/_01311_ ), .ZN(\mreg/_03932_ ) );
NAND3_X1 \mreg/_07185_ ( .A1(\mreg/_01177_ ), .A2(\mreg/_04575_ ), .A3(\mreg/_01178_ ), .ZN(\mreg/_01312_ ) );
NAND3_X1 \mreg/_07186_ ( .A1(\mreg/_01180_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04671_ ), .ZN(\mreg/_01313_ ) );
NAND3_X1 \mreg/_07187_ ( .A1(\mreg/_01182_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04607_ ), .ZN(\mreg/_01314_ ) );
INV_X1 \mreg/_07188_ ( .A(\mreg/_00033_ ), .ZN(\mreg/_01315_ ) );
NAND3_X1 \mreg/_07189_ ( .A1(\mreg/_01184_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_01315_ ), .ZN(\mreg/_01316_ ) );
AND4_X1 \mreg/_07190_ ( .A1(\mreg/_01312_ ), .A2(\mreg/_01313_ ), .A3(\mreg/_01314_ ), .A4(\mreg/_01316_ ), .ZN(\mreg/_01317_ ) );
BUF_X4 \mreg/_07191_ ( .A(\mreg/_01089_ ), .Z(\mreg/_01318_ ) );
NAND4_X1 \mreg/_07192_ ( .A1(\mreg/_01318_ ), .A2(\mreg/_01161_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04511_ ), .ZN(\mreg/_01319_ ) );
INV_X1 \mreg/_07193_ ( .A(\mreg/_04543_ ), .ZN(\mreg/_01320_ ) );
OAI21_X1 \mreg/_07194_ ( .A(\mreg/_01319_ ), .B1(\mreg/_01191_ ), .B2(\mreg/_01320_ ), .ZN(\mreg/_01321_ ) );
AOI221_X1 \mreg/_07195_ ( .A(\mreg/_01321_ ), .B1(\mreg/_04479_ ), .B2(\mreg/_01196_ ), .C1(\mreg/_04447_ ), .C2(\mreg/_01198_ ), .ZN(\mreg/_01322_ ) );
BUF_X4 \mreg/_07196_ ( .A(\mreg/_01090_ ), .Z(\mreg/_01323_ ) );
NAND3_X1 \mreg/_07197_ ( .A1(\mreg/_01323_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04383_ ), .ZN(\mreg/_01324_ ) );
NAND3_X1 \mreg/_07198_ ( .A1(\mreg/_01097_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04415_ ), .ZN(\mreg/_01325_ ) );
NAND2_X1 \mreg/_07199_ ( .A1(\mreg/_01324_ ), .A2(\mreg/_01325_ ), .ZN(\mreg/_01326_ ) );
AOI221_X1 \mreg/_07200_ ( .A(\mreg/_01326_ ), .B1(\mreg/_04351_ ), .B2(\mreg/_01205_ ), .C1(\mreg/_04319_ ), .C2(\mreg/_01207_ ), .ZN(\mreg/_01327_ ) );
NAND4_X1 \mreg/_07201_ ( .A1(\mreg/_01188_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04223_ ), .A4(\mreg/_01209_ ), .ZN(\mreg/_01328_ ) );
NAND4_X1 \mreg/_07202_ ( .A1(\mreg/_01211_ ), .A2(\mreg/_01212_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04255_ ), .ZN(\mreg/_01329_ ) );
NAND2_X1 \mreg/_07203_ ( .A1(\mreg/_01328_ ), .A2(\mreg/_01329_ ), .ZN(\mreg/_01330_ ) );
AOI221_X4 \mreg/_07204_ ( .A(\mreg/_01330_ ), .B1(\mreg/_01079_ ), .B2(\mreg/_04159_ ), .C1(\mreg/_04191_ ), .C2(\mreg/_01075_ ), .ZN(\mreg/_01331_ ) );
AND4_X1 \mreg/_07205_ ( .A1(\mreg/_01317_ ), .A2(\mreg/_01322_ ), .A3(\mreg/_01327_ ), .A4(\mreg/_01331_ ), .ZN(\mreg/_01332_ ) );
AND3_X1 \mreg/_07206_ ( .A1(\mreg/_01107_ ), .A2(\mreg/_01217_ ), .A3(\mreg/_04287_ ), .ZN(\mreg/_01333_ ) );
AOI221_X4 \mreg/_07207_ ( .A(\mreg/_01333_ ), .B1(\mreg/_01219_ ), .B2(\mreg/_04735_ ), .C1(\mreg/_04639_ ), .C2(\mreg/_01222_ ), .ZN(\mreg/_01334_ ) );
NAND3_X1 \mreg/_07208_ ( .A1(\mreg/_01059_ ), .A2(\mreg/_01287_ ), .A3(\mreg/_04799_ ), .ZN(\mreg/_01335_ ) );
NAND3_X1 \mreg/_07209_ ( .A1(\mreg/_01275_ ), .A2(\mreg/_01289_ ), .A3(\mreg/_04831_ ), .ZN(\mreg/_01336_ ) );
NAND3_X1 \mreg/_07210_ ( .A1(\mreg/_01281_ ), .A2(\mreg/_01306_ ), .A3(\mreg/_04863_ ), .ZN(\mreg/_01337_ ) );
BUF_X4 \mreg/_07211_ ( .A(\mreg/_01125_ ), .Z(\mreg/_01338_ ) );
BUF_X4 \mreg/_07212_ ( .A(\mreg/_01338_ ), .Z(\mreg/_01339_ ) );
NAND3_X1 \mreg/_07213_ ( .A1(\mreg/_01339_ ), .A2(\mreg/_01087_ ), .A3(\mreg/_04767_ ), .ZN(\mreg/_01340_ ) );
AND4_X1 \mreg/_07214_ ( .A1(\mreg/_01335_ ), .A2(\mreg/_01336_ ), .A3(\mreg/_01337_ ), .A4(\mreg/_01340_ ), .ZN(\mreg/_01341_ ) );
NAND3_X1 \mreg/_07215_ ( .A1(\mreg/_01158_ ), .A2(\mreg/_01233_ ), .A3(\mreg/_03967_ ), .ZN(\mreg/_01342_ ) );
NAND3_X1 \mreg/_07216_ ( .A1(\mreg/_01113_ ), .A2(\mreg/_01236_ ), .A3(\mreg/_03999_ ), .ZN(\mreg/_01343_ ) );
NAND3_X1 \mreg/_07217_ ( .A1(\mreg/_01155_ ), .A2(\mreg/_01239_ ), .A3(\mreg/_04927_ ), .ZN(\mreg/_01344_ ) );
NAND3_X1 \mreg/_07218_ ( .A1(\mreg/_01241_ ), .A2(\mreg/_01163_ ), .A3(\mreg/_04895_ ), .ZN(\mreg/_01345_ ) );
NAND4_X1 \mreg/_07219_ ( .A1(\mreg/_01342_ ), .A2(\mreg/_01343_ ), .A3(\mreg/_01344_ ), .A4(\mreg/_01345_ ), .ZN(\mreg/_01346_ ) );
NAND3_X1 \mreg/_07220_ ( .A1(\mreg/_01232_ ), .A2(\mreg/_01236_ ), .A3(\mreg/_04095_ ), .ZN(\mreg/_01347_ ) );
NAND3_X1 \mreg/_07221_ ( .A1(\mreg/_01238_ ), .A2(\mreg/_01236_ ), .A3(\mreg/_04127_ ), .ZN(\mreg/_01348_ ) );
NAND2_X1 \mreg/_07222_ ( .A1(\mreg/_01347_ ), .A2(\mreg/_01348_ ), .ZN(\mreg/_01349_ ) );
AND3_X1 \mreg/_07223_ ( .A1(\mreg/_01241_ ), .A2(\mreg/_04031_ ), .A3(\mreg/_01242_ ), .ZN(\mreg/_01350_ ) );
AND3_X1 \mreg/_07224_ ( .A1(\mreg/_01304_ ), .A2(\mreg/_01248_ ), .A3(\mreg/_04063_ ), .ZN(\mreg/_01351_ ) );
NOR4_X1 \mreg/_07225_ ( .A1(\mreg/_01346_ ), .A2(\mreg/_01349_ ), .A3(\mreg/_01350_ ), .A4(\mreg/_01351_ ), .ZN(\mreg/_01352_ ) );
NAND4_X1 \mreg/_07226_ ( .A1(\mreg/_01332_ ), .A2(\mreg/_01334_ ), .A3(\mreg/_01341_ ), .A4(\mreg/_01352_ ), .ZN(\mreg/_03935_ ) );
AND3_X1 \mreg/_07227_ ( .A1(\mreg/_01090_ ), .A2(\mreg/_01102_ ), .A3(\mreg/_04832_ ), .ZN(\mreg/_01353_ ) );
AND3_X1 \mreg/_07228_ ( .A1(\mreg/_01058_ ), .A2(\mreg/_01102_ ), .A3(\mreg/_04800_ ), .ZN(\mreg/_01354_ ) );
OR2_X1 \mreg/_07229_ ( .A1(\mreg/_01353_ ), .A2(\mreg/_01354_ ), .ZN(\mreg/_01355_ ) );
AOI221_X1 \mreg/_07230_ ( .A(\mreg/_01355_ ), .B1(\mreg/_04768_ ), .B2(\mreg/_01229_ ), .C1(\mreg/_04736_ ), .C2(\mreg/_01219_ ), .ZN(\mreg/_01356_ ) );
BUF_X2 \mreg/_07231_ ( .A(\mreg/_01102_ ), .Z(\mreg/_01357_ ) );
NAND3_X1 \mreg/_07232_ ( .A1(\mreg/_01146_ ), .A2(\mreg/_01357_ ), .A3(\mreg/_04064_ ), .ZN(\mreg/_01358_ ) );
NAND3_X1 \mreg/_07233_ ( .A1(\mreg/_01139_ ), .A2(\mreg/_01357_ ), .A3(\mreg/_04128_ ), .ZN(\mreg/_01359_ ) );
NAND2_X1 \mreg/_07234_ ( .A1(\mreg/_01358_ ), .A2(\mreg/_01359_ ), .ZN(\mreg/_01360_ ) );
AND2_X2 \mreg/_07235_ ( .A1(\mreg/_01117_ ), .A2(\mreg/_01108_ ), .ZN(\mreg/_01361_ ) );
AND2_X4 \mreg/_07236_ ( .A1(\mreg/_01121_ ), .A2(\mreg/_01108_ ), .ZN(\mreg/_01362_ ) );
BUF_X4 \mreg/_07237_ ( .A(\mreg/_01362_ ), .Z(\mreg/_01363_ ) );
AOI221_X1 \mreg/_07238_ ( .A(\mreg/_01360_ ), .B1(\mreg/_03968_ ), .B2(\mreg/_01361_ ), .C1(\mreg/_04928_ ), .C2(\mreg/_01363_ ), .ZN(\mreg/_01364_ ) );
BUF_X4 \mreg/_07239_ ( .A(\mreg/_01089_ ), .Z(\mreg/_01365_ ) );
BUF_X4 \mreg/_07240_ ( .A(\mreg/_01116_ ), .Z(\mreg/_01366_ ) );
NAND4_X1 \mreg/_07241_ ( .A1(\mreg/_01365_ ), .A2(\mreg/_01366_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04512_ ), .ZN(\mreg/_01367_ ) );
INV_X1 \mreg/_07242_ ( .A(\mreg/_04544_ ), .ZN(\mreg/_01368_ ) );
OAI21_X1 \mreg/_07243_ ( .A(\mreg/_01367_ ), .B1(\mreg/_01190_ ), .B2(\mreg/_01368_ ), .ZN(\mreg/_01369_ ) );
INV_X1 \mreg/_07244_ ( .A(\mreg/_00034_ ), .ZN(\mreg/_01370_ ) );
AOI221_X1 \mreg/_07245_ ( .A(\mreg/_01369_ ), .B1(\mreg/_01370_ ), .B2(\mreg/_01172_ ), .C1(\mreg/_04672_ ), .C2(\mreg/_01174_ ), .ZN(\mreg/_01371_ ) );
BUF_X4 \mreg/_07246_ ( .A(\mreg/_01062_ ), .Z(\mreg/_01372_ ) );
NAND4_X1 \mreg/_07247_ ( .A1(\mreg/_01365_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04224_ ), .A4(\mreg/_01372_ ), .ZN(\mreg/_01373_ ) );
BUF_X4 \mreg/_07248_ ( .A(\mreg/_01068_ ), .Z(\mreg/_01374_ ) );
INV_X1 \mreg/_07249_ ( .A(\mreg/_04256_ ), .ZN(\mreg/_01375_ ) );
OAI21_X1 \mreg/_07250_ ( .A(\mreg/_01373_ ), .B1(\mreg/_01374_ ), .B2(\mreg/_01375_ ), .ZN(\mreg/_01376_ ) );
BUF_X4 \mreg/_07251_ ( .A(\mreg/_01206_ ), .Z(\mreg/_01377_ ) );
AOI221_X1 \mreg/_07252_ ( .A(\mreg/_01376_ ), .B1(\mreg/_04352_ ), .B2(\mreg/_01204_ ), .C1(\mreg/_04320_ ), .C2(\mreg/_01377_ ), .ZN(\mreg/_01378_ ) );
NAND4_X1 \mreg/_07253_ ( .A1(\mreg/_01356_ ), .A2(\mreg/_01364_ ), .A3(\mreg/_01371_ ), .A4(\mreg/_01378_ ), .ZN(\mreg/_01379_ ) );
BUF_X2 \mreg/_07254_ ( .A(\mreg/_01097_ ), .Z(\mreg/_01380_ ) );
BUF_X2 \mreg/_07255_ ( .A(\mreg/_01380_ ), .Z(\mreg/_01381_ ) );
NAND3_X1 \mreg/_07256_ ( .A1(\mreg/_01381_ ), .A2(\mreg/_01239_ ), .A3(\mreg/_04864_ ), .ZN(\mreg/_01382_ ) );
BUF_X4 \mreg/_07257_ ( .A(\mreg/_01107_ ), .Z(\mreg/_01383_ ) );
BUF_X2 \mreg/_07258_ ( .A(\mreg/_01118_ ), .Z(\mreg/_01384_ ) );
NAND3_X1 \mreg/_07259_ ( .A1(\mreg/_01383_ ), .A2(\mreg/_01384_ ), .A3(\mreg/_04288_ ), .ZN(\mreg/_01385_ ) );
BUF_X4 \mreg/_07260_ ( .A(\mreg/_01064_ ), .Z(\mreg/_01386_ ) );
BUF_X2 \mreg/_07261_ ( .A(\mreg/_01122_ ), .Z(\mreg/_01387_ ) );
NAND3_X1 \mreg/_07262_ ( .A1(\mreg/_01386_ ), .A2(\mreg/_01387_ ), .A3(\mreg/_04640_ ), .ZN(\mreg/_01388_ ) );
NAND3_X1 \mreg/_07263_ ( .A1(\mreg/_01241_ ), .A2(\mreg/_01163_ ), .A3(\mreg/_04896_ ), .ZN(\mreg/_01389_ ) );
NAND4_X1 \mreg/_07264_ ( .A1(\mreg/_01382_ ), .A2(\mreg/_01385_ ), .A3(\mreg/_01388_ ), .A4(\mreg/_01389_ ), .ZN(\mreg/_01390_ ) );
BUF_X2 \mreg/_07265_ ( .A(\mreg/_01150_ ), .Z(\mreg/_01391_ ) );
NAND3_X1 \mreg/_07266_ ( .A1(\mreg/_01291_ ), .A2(\mreg/_04032_ ), .A3(\mreg/_01391_ ), .ZN(\mreg/_01392_ ) );
NAND2_X1 \mreg/_07267_ ( .A1(\mreg/_01142_ ), .A2(\mreg/_01118_ ), .ZN(\mreg/_01393_ ) );
INV_X1 \mreg/_07268_ ( .A(\mreg/_04096_ ), .ZN(\mreg/_01394_ ) );
INV_X1 \mreg/_07269_ ( .A(\mreg/_04000_ ), .ZN(\mreg/_01395_ ) );
NAND2_X2 \mreg/_07270_ ( .A1(\mreg/_01112_ ), .A2(\mreg/_01108_ ), .ZN(\mreg/_01396_ ) );
OAI221_X1 \mreg/_07271_ ( .A(\mreg/_01392_ ), .B1(\mreg/_01393_ ), .B2(\mreg/_01394_ ), .C1(\mreg/_01395_ ), .C2(\mreg/_01396_ ), .ZN(\mreg/_01397_ ) );
BUF_X8 \mreg/_07272_ ( .A(\mreg/_01090_ ), .Z(\mreg/_01398_ ) );
NAND3_X1 \mreg/_07273_ ( .A1(\mreg/_01398_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04384_ ), .ZN(\mreg/_01399_ ) );
NAND3_X1 \mreg/_07274_ ( .A1(\mreg/_01096_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04416_ ), .ZN(\mreg/_01400_ ) );
NAND2_X1 \mreg/_07275_ ( .A1(\mreg/_01399_ ), .A2(\mreg/_01400_ ), .ZN(\mreg/_01401_ ) );
AOI221_X1 \mreg/_07276_ ( .A(\mreg/_01401_ ), .B1(\mreg/_04192_ ), .B2(\mreg/_01074_ ), .C1(\mreg/_04160_ ), .C2(\mreg/_01079_ ), .ZN(\mreg/_01402_ ) );
AND3_X1 \mreg/_07277_ ( .A1(\mreg/_01255_ ), .A2(\mreg/_04448_ ), .A3(\mreg/_01127_ ), .ZN(\mreg/_01403_ ) );
AOI21_X1 \mreg/_07278_ ( .A(\mreg/_01403_ ), .B1(\mreg/_01196_ ), .B2(\mreg/_04480_ ), .ZN(\mreg/_01404_ ) );
NAND3_X1 \mreg/_07279_ ( .A1(\mreg/_01177_ ), .A2(\mreg/_04576_ ), .A3(\mreg/_01178_ ), .ZN(\mreg/_01405_ ) );
NAND3_X1 \mreg/_07280_ ( .A1(\mreg/_01304_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04608_ ), .ZN(\mreg/_01406_ ) );
NAND4_X1 \mreg/_07281_ ( .A1(\mreg/_01402_ ), .A2(\mreg/_01404_ ), .A3(\mreg/_01405_ ), .A4(\mreg/_01406_ ), .ZN(\mreg/_01407_ ) );
OR4_X1 \mreg/_07282_ ( .A1(\mreg/_01379_ ), .A2(\mreg/_01390_ ), .A3(\mreg/_01397_ ), .A4(\mreg/_01407_ ), .ZN(\mreg/_03936_ ) );
NAND3_X1 \mreg/_07283_ ( .A1(\mreg/_01084_ ), .A2(\mreg/_04577_ ), .A3(\mreg/_01299_ ), .ZN(\mreg/_01408_ ) );
NAND4_X1 \mreg/_07284_ ( .A1(\mreg/_01318_ ), .A2(\mreg/_01161_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04513_ ), .ZN(\mreg/_01409_ ) );
INV_X1 \mreg/_07285_ ( .A(\mreg/_04545_ ), .ZN(\mreg/_01410_ ) );
OAI21_X1 \mreg/_07286_ ( .A(\mreg/_01409_ ), .B1(\mreg/_01191_ ), .B2(\mreg/_01410_ ), .ZN(\mreg/_01411_ ) );
BUF_X4 \mreg/_07287_ ( .A(\mreg/_01195_ ), .Z(\mreg/_01412_ ) );
AOI221_X4 \mreg/_07288_ ( .A(\mreg/_01411_ ), .B1(\mreg/_04481_ ), .B2(\mreg/_01412_ ), .C1(\mreg/_04449_ ), .C2(\mreg/_01198_ ), .ZN(\mreg/_01413_ ) );
NAND3_X1 \mreg/_07289_ ( .A1(\mreg/_01305_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04609_ ), .ZN(\mreg/_01414_ ) );
AND3_X1 \mreg/_07290_ ( .A1(\mreg/_01143_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04673_ ), .ZN(\mreg/_01415_ ) );
INV_X1 \mreg/_07291_ ( .A(\mreg/_00035_ ), .ZN(\mreg/_01416_ ) );
AOI21_X1 \mreg/_07292_ ( .A(\mreg/_01415_ ), .B1(\mreg/_01416_ ), .B2(\mreg/_01173_ ), .ZN(\mreg/_01417_ ) );
AND4_X4 \mreg/_07293_ ( .A1(\mreg/_01408_ ), .A2(\mreg/_01413_ ), .A3(\mreg/_01414_ ), .A4(\mreg/_01417_ ), .ZN(\mreg/_01418_ ) );
NAND3_X1 \mreg/_07294_ ( .A1(\mreg/_01275_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04385_ ), .ZN(\mreg/_01419_ ) );
NAND4_X1 \mreg/_07295_ ( .A1(\mreg/_01365_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04225_ ), .A4(\mreg/_01372_ ), .ZN(\mreg/_01420_ ) );
INV_X1 \mreg/_07296_ ( .A(\mreg/_04257_ ), .ZN(\mreg/_01421_ ) );
OAI21_X1 \mreg/_07297_ ( .A(\mreg/_01420_ ), .B1(\mreg/_01374_ ), .B2(\mreg/_01421_ ), .ZN(\mreg/_01422_ ) );
AOI221_X4 \mreg/_07298_ ( .A(\mreg/_01422_ ), .B1(\mreg/_04193_ ), .B2(\mreg/_01074_ ), .C1(\mreg/_04161_ ), .C2(\mreg/_01079_ ), .ZN(\mreg/_01423_ ) );
NAND3_X1 \mreg/_07299_ ( .A1(\mreg/_01281_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04417_ ), .ZN(\mreg/_01424_ ) );
AND3_X1 \mreg/_07300_ ( .A1(\mreg/_01058_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04353_ ), .ZN(\mreg/_01425_ ) );
AOI21_X1 \mreg/_07301_ ( .A(\mreg/_01425_ ), .B1(\mreg/_04321_ ), .B2(\mreg/_01207_ ), .ZN(\mreg/_01426_ ) );
AND4_X1 \mreg/_07302_ ( .A1(\mreg/_01419_ ), .A2(\mreg/_01423_ ), .A3(\mreg/_01424_ ), .A4(\mreg/_01426_ ), .ZN(\mreg/_01427_ ) );
NAND3_X1 \mreg/_07303_ ( .A1(\mreg/_01383_ ), .A2(\mreg/_01287_ ), .A3(\mreg/_04289_ ), .ZN(\mreg/_01428_ ) );
AND3_X1 \mreg/_07304_ ( .A1(\mreg/_01098_ ), .A2(\mreg/_01133_ ), .A3(\mreg/_04865_ ), .ZN(\mreg/_01429_ ) );
AND2_X2 \mreg/_07305_ ( .A1(\mreg/_01090_ ), .A2(\mreg/_01102_ ), .ZN(\mreg/_01430_ ) );
BUF_X4 \mreg/_07306_ ( .A(\mreg/_01430_ ), .Z(\mreg/_01431_ ) );
AOI21_X1 \mreg/_07307_ ( .A(\mreg/_01429_ ), .B1(\mreg/_04833_ ), .B2(\mreg/_01431_ ), .ZN(\mreg/_01432_ ) );
AOI22_X1 \mreg/_07308_ ( .A1(\mreg/_04641_ ), .A2(\mreg/_01222_ ), .B1(\mreg/_01219_ ), .B2(\mreg/_04737_ ), .ZN(\mreg/_01433_ ) );
AOI22_X1 \mreg/_07309_ ( .A1(\mreg/_01228_ ), .A2(\mreg/_04801_ ), .B1(\mreg/_04769_ ), .B2(\mreg/_01229_ ), .ZN(\mreg/_01434_ ) );
AND4_X1 \mreg/_07310_ ( .A1(\mreg/_01428_ ), .A2(\mreg/_01432_ ), .A3(\mreg/_01433_ ), .A4(\mreg/_01434_ ), .ZN(\mreg/_01435_ ) );
BUF_X4 \mreg/_07311_ ( .A(\mreg/_01276_ ), .Z(\mreg/_01436_ ) );
NAND3_X1 \mreg/_07312_ ( .A1(\mreg/_01159_ ), .A2(\mreg/_01436_ ), .A3(\mreg/_03969_ ), .ZN(\mreg/_01437_ ) );
NAND3_X1 \mreg/_07313_ ( .A1(\mreg/_01338_ ), .A2(\mreg/_04033_ ), .A3(\mreg/_01151_ ), .ZN(\mreg/_01438_ ) );
NAND3_X1 \mreg/_07314_ ( .A1(\mreg/_01143_ ), .A2(\mreg/_01144_ ), .A3(\mreg/_04097_ ), .ZN(\mreg/_01439_ ) );
NAND3_X1 \mreg/_07315_ ( .A1(\mreg/_01148_ ), .A2(\mreg/_01133_ ), .A3(\mreg/_04065_ ), .ZN(\mreg/_01440_ ) );
NAND3_X1 \mreg/_07316_ ( .A1(\mreg/_01140_ ), .A2(\mreg/_01217_ ), .A3(\mreg/_04129_ ), .ZN(\mreg/_01441_ ) );
AND4_X1 \mreg/_07317_ ( .A1(\mreg/_01438_ ), .A2(\mreg/_01439_ ), .A3(\mreg/_01440_ ), .A4(\mreg/_01441_ ), .ZN(\mreg/_01442_ ) );
NAND3_X1 \mreg/_07318_ ( .A1(\mreg/_01165_ ), .A2(\mreg/_01306_ ), .A3(\mreg/_04001_ ), .ZN(\mreg/_01443_ ) );
AND3_X1 \mreg/_07319_ ( .A1(\mreg/_01126_ ), .A2(\mreg/_04897_ ), .A3(\mreg/_01162_ ), .ZN(\mreg/_01444_ ) );
AOI21_X1 \mreg/_07320_ ( .A(\mreg/_01444_ ), .B1(\mreg/_01363_ ), .B2(\mreg/_04929_ ), .ZN(\mreg/_01445_ ) );
AND4_X1 \mreg/_07321_ ( .A1(\mreg/_01437_ ), .A2(\mreg/_01442_ ), .A3(\mreg/_01443_ ), .A4(\mreg/_01445_ ), .ZN(\mreg/_01446_ ) );
NAND4_X1 \mreg/_07322_ ( .A1(\mreg/_01418_ ), .A2(\mreg/_01427_ ), .A3(\mreg/_01435_ ), .A4(\mreg/_01446_ ), .ZN(\mreg/_03937_ ) );
NAND3_X1 \mreg/_07323_ ( .A1(\mreg/_01177_ ), .A2(\mreg/_04578_ ), .A3(\mreg/_01178_ ), .ZN(\mreg/_01447_ ) );
NAND3_X1 \mreg/_07324_ ( .A1(\mreg/_01180_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04674_ ), .ZN(\mreg/_01448_ ) );
NAND3_X1 \mreg/_07325_ ( .A1(\mreg/_01182_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04610_ ), .ZN(\mreg/_01449_ ) );
INV_X1 \mreg/_07326_ ( .A(\mreg/_00036_ ), .ZN(\mreg/_01450_ ) );
NAND3_X1 \mreg/_07327_ ( .A1(\mreg/_01184_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_01450_ ), .ZN(\mreg/_01451_ ) );
AND4_X1 \mreg/_07328_ ( .A1(\mreg/_01447_ ), .A2(\mreg/_01448_ ), .A3(\mreg/_01449_ ), .A4(\mreg/_01451_ ), .ZN(\mreg/_01452_ ) );
BUF_X4 \mreg/_07329_ ( .A(\mreg/_01116_ ), .Z(\mreg/_01453_ ) );
NAND4_X1 \mreg/_07330_ ( .A1(\mreg/_01318_ ), .A2(\mreg/_01453_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04514_ ), .ZN(\mreg/_01454_ ) );
INV_X1 \mreg/_07331_ ( .A(\mreg/_04546_ ), .ZN(\mreg/_01455_ ) );
OAI21_X1 \mreg/_07332_ ( .A(\mreg/_01454_ ), .B1(\mreg/_01191_ ), .B2(\mreg/_01455_ ), .ZN(\mreg/_01456_ ) );
AOI221_X4 \mreg/_07333_ ( .A(\mreg/_01456_ ), .B1(\mreg/_04482_ ), .B2(\mreg/_01412_ ), .C1(\mreg/_04450_ ), .C2(\mreg/_01198_ ), .ZN(\mreg/_01457_ ) );
NAND3_X1 \mreg/_07334_ ( .A1(\mreg/_01323_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04386_ ), .ZN(\mreg/_01458_ ) );
NAND3_X1 \mreg/_07335_ ( .A1(\mreg/_01097_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04418_ ), .ZN(\mreg/_01459_ ) );
NAND2_X1 \mreg/_07336_ ( .A1(\mreg/_01458_ ), .A2(\mreg/_01459_ ), .ZN(\mreg/_01460_ ) );
AOI221_X4 \mreg/_07337_ ( .A(\mreg/_01460_ ), .B1(\mreg/_04354_ ), .B2(\mreg/_01205_ ), .C1(\mreg/_04322_ ), .C2(\mreg/_01207_ ), .ZN(\mreg/_01461_ ) );
NAND4_X1 \mreg/_07338_ ( .A1(\mreg/_01269_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04226_ ), .A4(\mreg/_01209_ ), .ZN(\mreg/_01462_ ) );
INV_X1 \mreg/_07339_ ( .A(\mreg/_04258_ ), .ZN(\mreg/_01463_ ) );
OAI21_X1 \mreg/_07340_ ( .A(\mreg/_01462_ ), .B1(\mreg/_01069_ ), .B2(\mreg/_01463_ ), .ZN(\mreg/_01464_ ) );
BUF_X4 \mreg/_07341_ ( .A(\mreg/_01074_ ), .Z(\mreg/_01465_ ) );
AOI221_X4 \mreg/_07342_ ( .A(\mreg/_01464_ ), .B1(\mreg/_04194_ ), .B2(\mreg/_01465_ ), .C1(\mreg/_04162_ ), .C2(\mreg/_01080_ ), .ZN(\mreg/_01466_ ) );
AND4_X2 \mreg/_07343_ ( .A1(\mreg/_01452_ ), .A2(\mreg/_01457_ ), .A3(\mreg/_01461_ ), .A4(\mreg/_01466_ ), .ZN(\mreg/_01467_ ) );
NAND3_X1 \mreg/_07344_ ( .A1(\mreg/_01275_ ), .A2(\mreg/_01277_ ), .A3(\mreg/_04834_ ), .ZN(\mreg/_01468_ ) );
AND3_X1 \mreg/_07345_ ( .A1(\mreg/_01072_ ), .A2(\mreg/_01103_ ), .A3(\mreg/_04290_ ), .ZN(\mreg/_01469_ ) );
AOI221_X4 \mreg/_07346_ ( .A(\mreg/_01469_ ), .B1(\mreg/_01106_ ), .B2(\mreg/_04738_ ), .C1(\mreg/_04642_ ), .C2(\mreg/_01221_ ), .ZN(\mreg/_01470_ ) );
NAND3_X1 \mreg/_07347_ ( .A1(\mreg/_01281_ ), .A2(\mreg/_01282_ ), .A3(\mreg/_04866_ ), .ZN(\mreg/_01471_ ) );
AOI22_X1 \mreg/_07348_ ( .A1(\mreg/_01284_ ), .A2(\mreg/_04802_ ), .B1(\mreg/_04770_ ), .B2(\mreg/_01230_ ), .ZN(\mreg/_01472_ ) );
AND4_X1 \mreg/_07349_ ( .A1(\mreg/_01468_ ), .A2(\mreg/_01470_ ), .A3(\mreg/_01471_ ), .A4(\mreg/_01472_ ), .ZN(\mreg/_01473_ ) );
NAND3_X1 \mreg/_07350_ ( .A1(\mreg/_01156_ ), .A2(\mreg/_01287_ ), .A3(\mreg/_04930_ ), .ZN(\mreg/_01474_ ) );
NAND3_X1 \mreg/_07351_ ( .A1(\mreg/_01159_ ), .A2(\mreg/_01289_ ), .A3(\mreg/_03970_ ), .ZN(\mreg/_01475_ ) );
NAND3_X1 \mreg/_07352_ ( .A1(\mreg/_01292_ ), .A2(\mreg/_01293_ ), .A3(\mreg/_04898_ ), .ZN(\mreg/_01476_ ) );
BUF_X2 \mreg/_07353_ ( .A(\mreg/_01130_ ), .Z(\mreg/_01477_ ) );
NAND3_X1 \mreg/_07354_ ( .A1(\mreg/_01165_ ), .A2(\mreg/_01477_ ), .A3(\mreg/_04002_ ), .ZN(\mreg/_01478_ ) );
AND4_X1 \mreg/_07355_ ( .A1(\mreg/_01474_ ), .A2(\mreg/_01475_ ), .A3(\mreg/_01476_ ), .A4(\mreg/_01478_ ), .ZN(\mreg/_01479_ ) );
AND3_X1 \mreg/_07356_ ( .A1(\mreg/_01232_ ), .A2(\mreg/_01233_ ), .A3(\mreg/_04098_ ), .ZN(\mreg/_01480_ ) );
AND3_X1 \mreg/_07357_ ( .A1(\mreg/_01235_ ), .A2(\mreg/_01239_ ), .A3(\mreg/_04066_ ), .ZN(\mreg/_01481_ ) );
AND3_X1 \mreg/_07358_ ( .A1(\mreg/_01238_ ), .A2(\mreg/_01248_ ), .A3(\mreg/_04130_ ), .ZN(\mreg/_01482_ ) );
AND3_X1 \mreg/_07359_ ( .A1(\mreg/_01250_ ), .A2(\mreg/_04034_ ), .A3(\mreg/_01391_ ), .ZN(\mreg/_01483_ ) );
NOR4_X1 \mreg/_07360_ ( .A1(\mreg/_01480_ ), .A2(\mreg/_01481_ ), .A3(\mreg/_01482_ ), .A4(\mreg/_01483_ ), .ZN(\mreg/_01484_ ) );
NAND4_X1 \mreg/_07361_ ( .A1(\mreg/_01467_ ), .A2(\mreg/_01473_ ), .A3(\mreg/_01479_ ), .A4(\mreg/_01484_ ), .ZN(\mreg/_03938_ ) );
NAND3_X1 \mreg/_07362_ ( .A1(\mreg/_01177_ ), .A2(\mreg/_04579_ ), .A3(\mreg/_01178_ ), .ZN(\mreg/_01485_ ) );
NAND3_X1 \mreg/_07363_ ( .A1(\mreg/_01180_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04675_ ), .ZN(\mreg/_01486_ ) );
NAND3_X1 \mreg/_07364_ ( .A1(\mreg/_01182_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04611_ ), .ZN(\mreg/_01487_ ) );
INV_X1 \mreg/_07365_ ( .A(\mreg/_00037_ ), .ZN(\mreg/_01488_ ) );
NAND3_X1 \mreg/_07366_ ( .A1(\mreg/_01184_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_01488_ ), .ZN(\mreg/_01489_ ) );
AND4_X1 \mreg/_07367_ ( .A1(\mreg/_01485_ ), .A2(\mreg/_01486_ ), .A3(\mreg/_01487_ ), .A4(\mreg/_01489_ ), .ZN(\mreg/_01490_ ) );
NAND4_X1 \mreg/_07368_ ( .A1(\mreg/_01318_ ), .A2(\mreg/_01453_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04515_ ), .ZN(\mreg/_01491_ ) );
INV_X1 \mreg/_07369_ ( .A(\mreg/_04547_ ), .ZN(\mreg/_01492_ ) );
OAI21_X1 \mreg/_07370_ ( .A(\mreg/_01491_ ), .B1(\mreg/_01191_ ), .B2(\mreg/_01492_ ), .ZN(\mreg/_01493_ ) );
AOI221_X4 \mreg/_07371_ ( .A(\mreg/_01493_ ), .B1(\mreg/_04483_ ), .B2(\mreg/_01412_ ), .C1(\mreg/_04451_ ), .C2(\mreg/_01198_ ), .ZN(\mreg/_01494_ ) );
NAND3_X1 \mreg/_07372_ ( .A1(\mreg/_01323_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04387_ ), .ZN(\mreg/_01495_ ) );
BUF_X4 \mreg/_07373_ ( .A(\mreg/_01096_ ), .Z(\mreg/_01496_ ) );
NAND3_X1 \mreg/_07374_ ( .A1(\mreg/_01496_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04419_ ), .ZN(\mreg/_01497_ ) );
NAND2_X1 \mreg/_07375_ ( .A1(\mreg/_01495_ ), .A2(\mreg/_01497_ ), .ZN(\mreg/_01498_ ) );
BUF_X4 \mreg/_07376_ ( .A(\mreg/_01206_ ), .Z(\mreg/_01499_ ) );
AOI221_X1 \mreg/_07377_ ( .A(\mreg/_01498_ ), .B1(\mreg/_04355_ ), .B2(\mreg/_01205_ ), .C1(\mreg/_04323_ ), .C2(\mreg/_01499_ ), .ZN(\mreg/_01500_ ) );
BUF_X4 \mreg/_07378_ ( .A(\mreg/_01089_ ), .Z(\mreg/_01501_ ) );
NAND4_X1 \mreg/_07379_ ( .A1(\mreg/_01501_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04227_ ), .A4(\mreg/_01209_ ), .ZN(\mreg/_01502_ ) );
INV_X1 \mreg/_07380_ ( .A(\mreg/_04259_ ), .ZN(\mreg/_01503_ ) );
OAI21_X1 \mreg/_07381_ ( .A(\mreg/_01502_ ), .B1(\mreg/_01069_ ), .B2(\mreg/_01503_ ), .ZN(\mreg/_01504_ ) );
BUF_X4 \mreg/_07382_ ( .A(\mreg/_01079_ ), .Z(\mreg/_01505_ ) );
AOI221_X4 \mreg/_07383_ ( .A(\mreg/_01504_ ), .B1(\mreg/_04195_ ), .B2(\mreg/_01465_ ), .C1(\mreg/_04163_ ), .C2(\mreg/_01505_ ), .ZN(\mreg/_01506_ ) );
AND4_X4 \mreg/_07384_ ( .A1(\mreg/_01490_ ), .A2(\mreg/_01494_ ), .A3(\mreg/_01500_ ), .A4(\mreg/_01506_ ), .ZN(\mreg/_01507_ ) );
NAND3_X1 \mreg/_07385_ ( .A1(\mreg/_01383_ ), .A2(\mreg/_01277_ ), .A3(\mreg/_04291_ ), .ZN(\mreg/_01508_ ) );
AOI22_X1 \mreg/_07386_ ( .A1(\mreg/_04643_ ), .A2(\mreg/_01222_ ), .B1(\mreg/_01219_ ), .B2(\mreg/_04739_ ), .ZN(\mreg/_01509_ ) );
AND3_X1 \mreg/_07387_ ( .A1(\mreg/_01098_ ), .A2(\mreg/_01133_ ), .A3(\mreg/_04867_ ), .ZN(\mreg/_01510_ ) );
AOI21_X1 \mreg/_07388_ ( .A(\mreg/_01510_ ), .B1(\mreg/_04835_ ), .B2(\mreg/_01431_ ), .ZN(\mreg/_01511_ ) );
AOI22_X1 \mreg/_07389_ ( .A1(\mreg/_01284_ ), .A2(\mreg/_04803_ ), .B1(\mreg/_04771_ ), .B2(\mreg/_01230_ ), .ZN(\mreg/_01512_ ) );
AND4_X1 \mreg/_07390_ ( .A1(\mreg/_01508_ ), .A2(\mreg/_01509_ ), .A3(\mreg/_01511_ ), .A4(\mreg/_01512_ ), .ZN(\mreg/_01513_ ) );
AND3_X1 \mreg/_07391_ ( .A1(\mreg/_01126_ ), .A2(\mreg/_04899_ ), .A3(\mreg/_01162_ ), .ZN(\mreg/_01514_ ) );
NAND3_X1 \mreg/_07392_ ( .A1(\mreg/_01117_ ), .A2(\mreg/_01118_ ), .A3(\mreg/_03971_ ), .ZN(\mreg/_01515_ ) );
INV_X1 \mreg/_07393_ ( .A(\mreg/_04003_ ), .ZN(\mreg/_01516_ ) );
OAI21_X1 \mreg/_07394_ ( .A(\mreg/_01515_ ), .B1(\mreg/_01516_ ), .B2(\mreg/_01396_ ), .ZN(\mreg/_01517_ ) );
AOI211_X4 \mreg/_07395_ ( .A(\mreg/_01514_ ), .B(\mreg/_01517_ ), .C1(\mreg/_04931_ ), .C2(\mreg/_01363_ ), .ZN(\mreg/_01518_ ) );
NAND3_X1 \mreg/_07396_ ( .A1(\mreg/_01298_ ), .A2(\mreg/_04035_ ), .A3(\mreg/_01299_ ), .ZN(\mreg/_01519_ ) );
NAND3_X1 \mreg/_07397_ ( .A1(\mreg/_01301_ ), .A2(\mreg/_01302_ ), .A3(\mreg/_04099_ ), .ZN(\mreg/_01520_ ) );
NAND3_X1 \mreg/_07398_ ( .A1(\mreg/_01305_ ), .A2(\mreg/_01306_ ), .A3(\mreg/_04067_ ), .ZN(\mreg/_01521_ ) );
NAND3_X1 \mreg/_07399_ ( .A1(\mreg/_01308_ ), .A2(\mreg/_01309_ ), .A3(\mreg/_04131_ ), .ZN(\mreg/_01522_ ) );
AND4_X1 \mreg/_07400_ ( .A1(\mreg/_01519_ ), .A2(\mreg/_01520_ ), .A3(\mreg/_01521_ ), .A4(\mreg/_01522_ ), .ZN(\mreg/_01523_ ) );
NAND4_X1 \mreg/_07401_ ( .A1(\mreg/_01507_ ), .A2(\mreg/_01513_ ), .A3(\mreg/_01518_ ), .A4(\mreg/_01523_ ), .ZN(\mreg/_03939_ ) );
NAND3_X1 \mreg/_07402_ ( .A1(\mreg/_01067_ ), .A2(\mreg/_01109_ ), .A3(\mreg/_04740_ ), .ZN(\mreg/_01524_ ) );
NAND3_X1 \mreg/_07403_ ( .A1(\mreg/_01125_ ), .A2(\mreg/_01086_ ), .A3(\mreg/_04772_ ), .ZN(\mreg/_01525_ ) );
NAND2_X1 \mreg/_07404_ ( .A1(\mreg/_01524_ ), .A2(\mreg/_01525_ ), .ZN(\mreg/_01526_ ) );
AOI221_X4 \mreg/_07405_ ( .A(\mreg/_01526_ ), .B1(\mreg/_04836_ ), .B2(\mreg/_01431_ ), .C1(\mreg/_04804_ ), .C2(\mreg/_01228_ ), .ZN(\mreg/_01527_ ) );
NAND4_X1 \mreg/_07406_ ( .A1(\mreg/_01318_ ), .A2(\mreg/_01453_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04516_ ), .ZN(\mreg/_01528_ ) );
INV_X1 \mreg/_07407_ ( .A(\mreg/_04548_ ), .ZN(\mreg/_01529_ ) );
OAI21_X1 \mreg/_07408_ ( .A(\mreg/_01528_ ), .B1(\mreg/_01191_ ), .B2(\mreg/_01529_ ), .ZN(\mreg/_01530_ ) );
INV_X1 \mreg/_07409_ ( .A(\mreg/_00038_ ), .ZN(\mreg/_01531_ ) );
AOI221_X4 \mreg/_07410_ ( .A(\mreg/_01530_ ), .B1(\mreg/_01531_ ), .B2(\mreg/_01172_ ), .C1(\mreg/_04676_ ), .C2(\mreg/_01175_ ), .ZN(\mreg/_01532_ ) );
NAND3_X1 \mreg/_07411_ ( .A1(\mreg/_01146_ ), .A2(\mreg/_01103_ ), .A3(\mreg/_04068_ ), .ZN(\mreg/_01533_ ) );
NAND3_X1 \mreg/_07412_ ( .A1(\mreg/_01139_ ), .A2(\mreg/_01103_ ), .A3(\mreg/_04132_ ), .ZN(\mreg/_01534_ ) );
NAND2_X1 \mreg/_07413_ ( .A1(\mreg/_01533_ ), .A2(\mreg/_01534_ ), .ZN(\mreg/_01535_ ) );
AOI221_X4 \mreg/_07414_ ( .A(\mreg/_01535_ ), .B1(\mreg/_03972_ ), .B2(\mreg/_01361_ ), .C1(\mreg/_04932_ ), .C2(\mreg/_01363_ ), .ZN(\mreg/_01536_ ) );
NAND4_X1 \mreg/_07415_ ( .A1(\mreg/_01501_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04228_ ), .A4(\mreg/_01209_ ), .ZN(\mreg/_01537_ ) );
INV_X1 \mreg/_07416_ ( .A(\mreg/_04260_ ), .ZN(\mreg/_01538_ ) );
OAI21_X1 \mreg/_07417_ ( .A(\mreg/_01537_ ), .B1(\mreg/_01069_ ), .B2(\mreg/_01538_ ), .ZN(\mreg/_01539_ ) );
AOI221_X4 \mreg/_07418_ ( .A(\mreg/_01539_ ), .B1(\mreg/_04356_ ), .B2(\mreg/_01204_ ), .C1(\mreg/_04324_ ), .C2(\mreg/_01377_ ), .ZN(\mreg/_01540_ ) );
AND4_X4 \mreg/_07419_ ( .A1(\mreg/_01527_ ), .A2(\mreg/_01532_ ), .A3(\mreg/_01536_ ), .A4(\mreg/_01540_ ), .ZN(\mreg/_01541_ ) );
NAND3_X1 \mreg/_07420_ ( .A1(\mreg/_01339_ ), .A2(\mreg/_04036_ ), .A3(\mreg/_01242_ ), .ZN(\mreg/_01542_ ) );
INV_X1 \mreg/_07421_ ( .A(\mreg/_04100_ ), .ZN(\mreg/_01543_ ) );
INV_X1 \mreg/_07422_ ( .A(\mreg/_04004_ ), .ZN(\mreg/_01544_ ) );
OAI221_X1 \mreg/_07423_ ( .A(\mreg/_01542_ ), .B1(\mreg/_01393_ ), .B2(\mreg/_01543_ ), .C1(\mreg/_01544_ ), .C2(\mreg/_01396_ ), .ZN(\mreg/_01545_ ) );
AND3_X1 \mreg/_07424_ ( .A1(\mreg/_01381_ ), .A2(\mreg/_01233_ ), .A3(\mreg/_04868_ ), .ZN(\mreg/_01546_ ) );
AND3_X1 \mreg/_07425_ ( .A1(\mreg/_01241_ ), .A2(\mreg/_04900_ ), .A3(\mreg/_01163_ ), .ZN(\mreg/_01547_ ) );
NAND3_X1 \mreg/_07426_ ( .A1(\mreg/_01383_ ), .A2(\mreg/_01384_ ), .A3(\mreg/_04292_ ), .ZN(\mreg/_01548_ ) );
NAND3_X1 \mreg/_07427_ ( .A1(\mreg/_01386_ ), .A2(\mreg/_01387_ ), .A3(\mreg/_04644_ ), .ZN(\mreg/_01549_ ) );
NAND2_X1 \mreg/_07428_ ( .A1(\mreg/_01548_ ), .A2(\mreg/_01549_ ), .ZN(\mreg/_01550_ ) );
NOR4_X1 \mreg/_07429_ ( .A1(\mreg/_01545_ ), .A2(\mreg/_01546_ ), .A3(\mreg/_01547_ ), .A4(\mreg/_01550_ ), .ZN(\mreg/_01551_ ) );
NAND3_X1 \mreg/_07430_ ( .A1(\mreg/_01156_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04484_ ), .ZN(\mreg/_01552_ ) );
NAND3_X1 \mreg/_07431_ ( .A1(\mreg/_01305_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04612_ ), .ZN(\mreg/_01553_ ) );
NAND3_X1 \mreg/_07432_ ( .A1(\mreg/_01084_ ), .A2(\mreg/_04580_ ), .A3(\mreg/_01242_ ), .ZN(\mreg/_01554_ ) );
NAND3_X1 \mreg/_07433_ ( .A1(\mreg/_01084_ ), .A2(\mreg/_04452_ ), .A3(\mreg/_01163_ ), .ZN(\mreg/_01555_ ) );
AND4_X1 \mreg/_07434_ ( .A1(\mreg/_01552_ ), .A2(\mreg/_01553_ ), .A3(\mreg/_01554_ ), .A4(\mreg/_01555_ ), .ZN(\mreg/_01556_ ) );
NAND3_X1 \mreg/_07435_ ( .A1(\mreg/_01091_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04388_ ), .ZN(\mreg/_01557_ ) );
NAND3_X1 \mreg/_07436_ ( .A1(\mreg/_01380_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04420_ ), .ZN(\mreg/_01558_ ) );
NAND2_X1 \mreg/_07437_ ( .A1(\mreg/_01557_ ), .A2(\mreg/_01558_ ), .ZN(\mreg/_01559_ ) );
AOI221_X4 \mreg/_07438_ ( .A(\mreg/_01559_ ), .B1(\mreg/_04196_ ), .B2(\mreg/_01075_ ), .C1(\mreg/_04164_ ), .C2(\mreg/_01080_ ), .ZN(\mreg/_01560_ ) );
NAND4_X1 \mreg/_07439_ ( .A1(\mreg/_01541_ ), .A2(\mreg/_01551_ ), .A3(\mreg/_01556_ ), .A4(\mreg/_01560_ ), .ZN(\mreg/_03940_ ) );
AND3_X1 \mreg/_07440_ ( .A1(\mreg/_01090_ ), .A2(\mreg/_01102_ ), .A3(\mreg/_04837_ ), .ZN(\mreg/_01561_ ) );
AND3_X1 \mreg/_07441_ ( .A1(\mreg/_01058_ ), .A2(\mreg/_01102_ ), .A3(\mreg/_04805_ ), .ZN(\mreg/_01562_ ) );
OR2_X1 \mreg/_07442_ ( .A1(\mreg/_01561_ ), .A2(\mreg/_01562_ ), .ZN(\mreg/_01563_ ) );
AOI221_X4 \mreg/_07443_ ( .A(\mreg/_01563_ ), .B1(\mreg/_04773_ ), .B2(\mreg/_01229_ ), .C1(\mreg/_04741_ ), .C2(\mreg/_01106_ ), .ZN(\mreg/_01564_ ) );
NAND3_X1 \mreg/_07444_ ( .A1(\mreg/_01146_ ), .A2(\mreg/_01357_ ), .A3(\mreg/_04069_ ), .ZN(\mreg/_01565_ ) );
NAND3_X1 \mreg/_07445_ ( .A1(\mreg/_01139_ ), .A2(\mreg/_01357_ ), .A3(\mreg/_04133_ ), .ZN(\mreg/_01566_ ) );
NAND2_X1 \mreg/_07446_ ( .A1(\mreg/_01565_ ), .A2(\mreg/_01566_ ), .ZN(\mreg/_01567_ ) );
AOI221_X4 \mreg/_07447_ ( .A(\mreg/_01567_ ), .B1(\mreg/_03973_ ), .B2(\mreg/_01361_ ), .C1(\mreg/_04933_ ), .C2(\mreg/_01363_ ), .ZN(\mreg/_01568_ ) );
NAND4_X1 \mreg/_07448_ ( .A1(\mreg/_01365_ ), .A2(\mreg/_01366_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04517_ ), .ZN(\mreg/_01569_ ) );
INV_X1 \mreg/_07449_ ( .A(\mreg/_04549_ ), .ZN(\mreg/_01570_ ) );
OAI21_X1 \mreg/_07450_ ( .A(\mreg/_01569_ ), .B1(\mreg/_01190_ ), .B2(\mreg/_01570_ ), .ZN(\mreg/_01571_ ) );
INV_X1 \mreg/_07451_ ( .A(\mreg/_00039_ ), .ZN(\mreg/_01572_ ) );
AOI221_X1 \mreg/_07452_ ( .A(\mreg/_01571_ ), .B1(\mreg/_01572_ ), .B2(\mreg/_01172_ ), .C1(\mreg/_04677_ ), .C2(\mreg/_01174_ ), .ZN(\mreg/_01573_ ) );
NAND4_X1 \mreg/_07453_ ( .A1(\mreg/_01365_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04229_ ), .A4(\mreg/_01062_ ), .ZN(\mreg/_01574_ ) );
INV_X1 \mreg/_07454_ ( .A(\mreg/_04261_ ), .ZN(\mreg/_01575_ ) );
OAI21_X1 \mreg/_07455_ ( .A(\mreg/_01574_ ), .B1(\mreg/_01068_ ), .B2(\mreg/_01575_ ), .ZN(\mreg/_01576_ ) );
AOI221_X4 \mreg/_07456_ ( .A(\mreg/_01576_ ), .B1(\mreg/_04357_ ), .B2(\mreg/_01204_ ), .C1(\mreg/_04325_ ), .C2(\mreg/_01377_ ), .ZN(\mreg/_01577_ ) );
NAND4_X1 \mreg/_07457_ ( .A1(\mreg/_01564_ ), .A2(\mreg/_01568_ ), .A3(\mreg/_01573_ ), .A4(\mreg/_01577_ ), .ZN(\mreg/_01578_ ) );
NAND3_X1 \mreg/_07458_ ( .A1(\mreg/_01381_ ), .A2(\mreg/_01239_ ), .A3(\mreg/_04869_ ), .ZN(\mreg/_01579_ ) );
NAND3_X1 \mreg/_07459_ ( .A1(\mreg/_01383_ ), .A2(\mreg/_01384_ ), .A3(\mreg/_04293_ ), .ZN(\mreg/_01580_ ) );
NAND3_X1 \mreg/_07460_ ( .A1(\mreg/_01386_ ), .A2(\mreg/_01387_ ), .A3(\mreg/_04645_ ), .ZN(\mreg/_01581_ ) );
NAND3_X1 \mreg/_07461_ ( .A1(\mreg/_01241_ ), .A2(\mreg/_01163_ ), .A3(\mreg/_04901_ ), .ZN(\mreg/_01582_ ) );
NAND4_X1 \mreg/_07462_ ( .A1(\mreg/_01579_ ), .A2(\mreg/_01580_ ), .A3(\mreg/_01581_ ), .A4(\mreg/_01582_ ), .ZN(\mreg/_01583_ ) );
NAND3_X1 \mreg/_07463_ ( .A1(\mreg/_01232_ ), .A2(\mreg/_01276_ ), .A3(\mreg/_04101_ ), .ZN(\mreg/_01584_ ) );
NAND3_X1 \mreg/_07464_ ( .A1(\mreg/_01291_ ), .A2(\mreg/_04037_ ), .A3(\mreg/_01178_ ), .ZN(\mreg/_01585_ ) );
INV_X1 \mreg/_07465_ ( .A(\mreg/_04005_ ), .ZN(\mreg/_01586_ ) );
OAI211_X2 \mreg/_07466_ ( .A(\mreg/_01584_ ), .B(\mreg/_01585_ ), .C1(\mreg/_01396_ ), .C2(\mreg/_01586_ ), .ZN(\mreg/_01587_ ) );
NAND3_X1 \mreg/_07467_ ( .A1(\mreg/_01398_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04389_ ), .ZN(\mreg/_01588_ ) );
NAND3_X1 \mreg/_07468_ ( .A1(\mreg/_01096_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04421_ ), .ZN(\mreg/_01589_ ) );
NAND2_X1 \mreg/_07469_ ( .A1(\mreg/_01588_ ), .A2(\mreg/_01589_ ), .ZN(\mreg/_01590_ ) );
AOI221_X1 \mreg/_07470_ ( .A(\mreg/_01590_ ), .B1(\mreg/_04197_ ), .B2(\mreg/_01074_ ), .C1(\mreg/_04165_ ), .C2(\mreg/_01079_ ), .ZN(\mreg/_01591_ ) );
AND3_X1 \mreg/_07471_ ( .A1(\mreg/_01255_ ), .A2(\mreg/_04453_ ), .A3(\mreg/_01127_ ), .ZN(\mreg/_01592_ ) );
AOI21_X1 \mreg/_07472_ ( .A(\mreg/_01592_ ), .B1(\mreg/_01196_ ), .B2(\mreg/_04485_ ), .ZN(\mreg/_01593_ ) );
NAND3_X1 \mreg/_07473_ ( .A1(\mreg/_01177_ ), .A2(\mreg/_04581_ ), .A3(\mreg/_01178_ ), .ZN(\mreg/_01594_ ) );
NAND3_X1 \mreg/_07474_ ( .A1(\mreg/_01304_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04613_ ), .ZN(\mreg/_01595_ ) );
NAND4_X1 \mreg/_07475_ ( .A1(\mreg/_01591_ ), .A2(\mreg/_01593_ ), .A3(\mreg/_01594_ ), .A4(\mreg/_01595_ ), .ZN(\mreg/_01596_ ) );
OR4_X2 \mreg/_07476_ ( .A1(\mreg/_01578_ ), .A2(\mreg/_01583_ ), .A3(\mreg/_01587_ ), .A4(\mreg/_01596_ ), .ZN(\mreg/_03941_ ) );
BUF_X4 \mreg/_07477_ ( .A(\mreg/_01150_ ), .Z(\mreg/_01597_ ) );
NAND3_X1 \mreg/_07478_ ( .A1(\mreg/_01083_ ), .A2(\mreg/_04551_ ), .A3(\mreg/_01597_ ), .ZN(\mreg/_01598_ ) );
NAND3_X1 \mreg/_07479_ ( .A1(\mreg/_01180_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04647_ ), .ZN(\mreg/_01599_ ) );
NAND3_X1 \mreg/_07480_ ( .A1(\mreg/_01182_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04583_ ), .ZN(\mreg/_01600_ ) );
INV_X1 \mreg/_07481_ ( .A(\mreg/_00040_ ), .ZN(\mreg/_01601_ ) );
NAND3_X1 \mreg/_07482_ ( .A1(\mreg/_01184_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_01601_ ), .ZN(\mreg/_01602_ ) );
AND4_X1 \mreg/_07483_ ( .A1(\mreg/_01598_ ), .A2(\mreg/_01599_ ), .A3(\mreg/_01600_ ), .A4(\mreg/_01602_ ), .ZN(\mreg/_01603_ ) );
NAND4_X1 \mreg/_07484_ ( .A1(\mreg/_01318_ ), .A2(\mreg/_01453_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04487_ ), .ZN(\mreg/_01604_ ) );
INV_X1 \mreg/_07485_ ( .A(\mreg/_04519_ ), .ZN(\mreg/_01605_ ) );
OAI21_X1 \mreg/_07486_ ( .A(\mreg/_01604_ ), .B1(\mreg/_01191_ ), .B2(\mreg/_01605_ ), .ZN(\mreg/_01606_ ) );
AOI221_X4 \mreg/_07487_ ( .A(\mreg/_01606_ ), .B1(\mreg/_04455_ ), .B2(\mreg/_01412_ ), .C1(\mreg/_04423_ ), .C2(\mreg/_01198_ ), .ZN(\mreg/_01607_ ) );
NAND3_X1 \mreg/_07488_ ( .A1(\mreg/_01323_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04359_ ), .ZN(\mreg/_01608_ ) );
NAND3_X1 \mreg/_07489_ ( .A1(\mreg/_01496_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04391_ ), .ZN(\mreg/_01609_ ) );
NAND2_X1 \mreg/_07490_ ( .A1(\mreg/_01608_ ), .A2(\mreg/_01609_ ), .ZN(\mreg/_01610_ ) );
BUF_X4 \mreg/_07491_ ( .A(\mreg/_01203_ ), .Z(\mreg/_01611_ ) );
AOI221_X4 \mreg/_07492_ ( .A(\mreg/_01610_ ), .B1(\mreg/_04327_ ), .B2(\mreg/_01611_ ), .C1(\mreg/_04295_ ), .C2(\mreg/_01499_ ), .ZN(\mreg/_01612_ ) );
NAND4_X1 \mreg/_07493_ ( .A1(\mreg/_01501_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04199_ ), .A4(\mreg/_01209_ ), .ZN(\mreg/_01613_ ) );
INV_X1 \mreg/_07494_ ( .A(\mreg/_04231_ ), .ZN(\mreg/_01614_ ) );
OAI21_X1 \mreg/_07495_ ( .A(\mreg/_01613_ ), .B1(\mreg/_01069_ ), .B2(\mreg/_01614_ ), .ZN(\mreg/_01615_ ) );
AOI221_X4 \mreg/_07496_ ( .A(\mreg/_01615_ ), .B1(\mreg/_04167_ ), .B2(\mreg/_01465_ ), .C1(\mreg/_04135_ ), .C2(\mreg/_01505_ ), .ZN(\mreg/_01616_ ) );
AND4_X2 \mreg/_07497_ ( .A1(\mreg/_01603_ ), .A2(\mreg/_01607_ ), .A3(\mreg/_01612_ ), .A4(\mreg/_01616_ ), .ZN(\mreg/_01617_ ) );
NAND3_X1 \mreg/_07498_ ( .A1(\mreg/_01275_ ), .A2(\mreg/_01277_ ), .A3(\mreg/_04807_ ), .ZN(\mreg/_01618_ ) );
AOI22_X1 \mreg/_07499_ ( .A1(\mreg/_01284_ ), .A2(\mreg/_04775_ ), .B1(\mreg/_04743_ ), .B2(\mreg/_01230_ ), .ZN(\mreg/_01619_ ) );
NAND3_X1 \mreg/_07500_ ( .A1(\mreg/_01281_ ), .A2(\mreg/_01282_ ), .A3(\mreg/_04839_ ), .ZN(\mreg/_01620_ ) );
BUF_X4 \mreg/_07501_ ( .A(\mreg/_01107_ ), .Z(\mreg/_01621_ ) );
BUF_X2 \mreg/_07502_ ( .A(\mreg/_01109_ ), .Z(\mreg/_01622_ ) );
NAND3_X1 \mreg/_07503_ ( .A1(\mreg/_01621_ ), .A2(\mreg/_01622_ ), .A3(\mreg/_04263_ ), .ZN(\mreg/_01623_ ) );
NAND3_X1 \mreg/_07504_ ( .A1(\mreg/_01386_ ), .A2(\mreg/_01622_ ), .A3(\mreg/_04615_ ), .ZN(\mreg/_01624_ ) );
NAND3_X1 \mreg/_07505_ ( .A1(\mreg/_01067_ ), .A2(\mreg/_01130_ ), .A3(\mreg/_04711_ ), .ZN(\mreg/_01625_ ) );
AND3_X1 \mreg/_07506_ ( .A1(\mreg/_01623_ ), .A2(\mreg/_01624_ ), .A3(\mreg/_01625_ ), .ZN(\mreg/_01626_ ) );
AND4_X1 \mreg/_07507_ ( .A1(\mreg/_01618_ ), .A2(\mreg/_01619_ ), .A3(\mreg/_01620_ ), .A4(\mreg/_01626_ ), .ZN(\mreg/_01627_ ) );
AND3_X1 \mreg/_07508_ ( .A1(\mreg/_01113_ ), .A2(\mreg/_01477_ ), .A3(\mreg/_03975_ ), .ZN(\mreg/_01628_ ) );
AND3_X1 \mreg/_07509_ ( .A1(\mreg/_01158_ ), .A2(\mreg/_01236_ ), .A3(\mreg/_03943_ ), .ZN(\mreg/_01629_ ) );
AND3_X1 \mreg/_07510_ ( .A1(\mreg/_01155_ ), .A2(\mreg/_01387_ ), .A3(\mreg/_04903_ ), .ZN(\mreg/_01630_ ) );
AND3_X1 \mreg/_07511_ ( .A1(\mreg/_01250_ ), .A2(\mreg/_04871_ ), .A3(\mreg/_01251_ ), .ZN(\mreg/_01631_ ) );
NOR4_X1 \mreg/_07512_ ( .A1(\mreg/_01628_ ), .A2(\mreg/_01629_ ), .A3(\mreg/_01630_ ), .A4(\mreg/_01631_ ), .ZN(\mreg/_01632_ ) );
AND3_X1 \mreg/_07513_ ( .A1(\mreg/_01232_ ), .A2(\mreg/_01233_ ), .A3(\mreg/_04071_ ), .ZN(\mreg/_01633_ ) );
AND3_X1 \mreg/_07514_ ( .A1(\mreg/_01235_ ), .A2(\mreg/_01384_ ), .A3(\mreg/_04039_ ), .ZN(\mreg/_01634_ ) );
AND3_X1 \mreg/_07515_ ( .A1(\mreg/_01238_ ), .A2(\mreg/_01248_ ), .A3(\mreg/_04103_ ), .ZN(\mreg/_01635_ ) );
AND3_X1 \mreg/_07516_ ( .A1(\mreg/_01250_ ), .A2(\mreg/_04007_ ), .A3(\mreg/_01391_ ), .ZN(\mreg/_01636_ ) );
NOR4_X1 \mreg/_07517_ ( .A1(\mreg/_01633_ ), .A2(\mreg/_01634_ ), .A3(\mreg/_01635_ ), .A4(\mreg/_01636_ ), .ZN(\mreg/_01637_ ) );
NAND4_X1 \mreg/_07518_ ( .A1(\mreg/_01617_ ), .A2(\mreg/_01627_ ), .A3(\mreg/_01632_ ), .A4(\mreg/_01637_ ), .ZN(\mreg/_03911_ ) );
AND3_X1 \mreg/_07519_ ( .A1(\mreg/_01107_ ), .A2(\mreg/_01109_ ), .A3(\mreg/_04264_ ), .ZN(\mreg/_01638_ ) );
AOI221_X4 \mreg/_07520_ ( .A(\mreg/_01638_ ), .B1(\mreg/_01106_ ), .B2(\mreg/_04712_ ), .C1(\mreg/_04616_ ), .C2(\mreg/_01222_ ), .ZN(\mreg/_01639_ ) );
NAND3_X1 \mreg/_07521_ ( .A1(\mreg/_01121_ ), .A2(\mreg/_01276_ ), .A3(\mreg/_04904_ ), .ZN(\mreg/_01640_ ) );
NAND3_X1 \mreg/_07522_ ( .A1(\mreg/_01158_ ), .A2(\mreg/_01622_ ), .A3(\mreg/_03944_ ), .ZN(\mreg/_01641_ ) );
NAND3_X1 \mreg/_07523_ ( .A1(\mreg/_01338_ ), .A2(\mreg/_01251_ ), .A3(\mreg/_04872_ ), .ZN(\mreg/_01642_ ) );
NAND3_X1 \mreg/_07524_ ( .A1(\mreg/_01113_ ), .A2(\mreg/_01114_ ), .A3(\mreg/_03976_ ), .ZN(\mreg/_01643_ ) );
AND4_X1 \mreg/_07525_ ( .A1(\mreg/_01640_ ), .A2(\mreg/_01641_ ), .A3(\mreg/_01642_ ), .A4(\mreg/_01643_ ), .ZN(\mreg/_01644_ ) );
NAND3_X1 \mreg/_07526_ ( .A1(\mreg/_01059_ ), .A2(\mreg/_01622_ ), .A3(\mreg/_04776_ ), .ZN(\mreg/_01645_ ) );
NAND3_X1 \mreg/_07527_ ( .A1(\mreg/_01092_ ), .A2(\mreg/_01130_ ), .A3(\mreg/_04808_ ), .ZN(\mreg/_01646_ ) );
NAND3_X1 \mreg/_07528_ ( .A1(\mreg/_01098_ ), .A2(\mreg/_01114_ ), .A3(\mreg/_04840_ ), .ZN(\mreg/_01647_ ) );
NAND3_X1 \mreg/_07529_ ( .A1(\mreg/_01338_ ), .A2(\mreg/_01086_ ), .A3(\mreg/_04744_ ), .ZN(\mreg/_01648_ ) );
AND4_X1 \mreg/_07530_ ( .A1(\mreg/_01645_ ), .A2(\mreg/_01646_ ), .A3(\mreg/_01647_ ), .A4(\mreg/_01648_ ), .ZN(\mreg/_01649_ ) );
NAND3_X1 \mreg/_07531_ ( .A1(\mreg/_01291_ ), .A2(\mreg/_04008_ ), .A3(\mreg/_01597_ ), .ZN(\mreg/_01650_ ) );
NAND3_X1 \mreg/_07532_ ( .A1(\mreg/_01143_ ), .A2(\mreg/_01114_ ), .A3(\mreg/_04072_ ), .ZN(\mreg/_01651_ ) );
NAND3_X1 \mreg/_07533_ ( .A1(\mreg/_01148_ ), .A2(\mreg/_01114_ ), .A3(\mreg/_04040_ ), .ZN(\mreg/_01652_ ) );
NAND3_X1 \mreg/_07534_ ( .A1(\mreg/_01140_ ), .A2(\mreg/_01144_ ), .A3(\mreg/_04104_ ), .ZN(\mreg/_01653_ ) );
AND4_X1 \mreg/_07535_ ( .A1(\mreg/_01650_ ), .A2(\mreg/_01651_ ), .A3(\mreg/_01652_ ), .A4(\mreg/_01653_ ), .ZN(\mreg/_01654_ ) );
AND4_X1 \mreg/_07536_ ( .A1(\mreg/_01639_ ), .A2(\mreg/_01644_ ), .A3(\mreg/_01649_ ), .A4(\mreg/_01654_ ), .ZN(\mreg/_01655_ ) );
NAND3_X1 \mreg/_07537_ ( .A1(\mreg/_01084_ ), .A2(\mreg/_04552_ ), .A3(\mreg/_01299_ ), .ZN(\mreg/_01656_ ) );
NAND4_X1 \mreg/_07538_ ( .A1(\mreg/_01188_ ), .A2(\mreg/_01161_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04488_ ), .ZN(\mreg/_01657_ ) );
NAND4_X1 \mreg/_07539_ ( .A1(\mreg/_01161_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_01066_ ), .A4(\mreg/_04520_ ), .ZN(\mreg/_01658_ ) );
NAND2_X1 \mreg/_07540_ ( .A1(\mreg/_01657_ ), .A2(\mreg/_01658_ ), .ZN(\mreg/_01659_ ) );
BUF_X4 \mreg/_07541_ ( .A(\mreg/_01197_ ), .Z(\mreg/_01660_ ) );
AOI221_X4 \mreg/_07542_ ( .A(\mreg/_01659_ ), .B1(\mreg/_01660_ ), .B2(\mreg/_04424_ ), .C1(\mreg/_04456_ ), .C2(\mreg/_01196_ ), .ZN(\mreg/_01661_ ) );
NAND3_X1 \mreg/_07543_ ( .A1(\mreg/_01305_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04584_ ), .ZN(\mreg/_01662_ ) );
AND3_X1 \mreg/_07544_ ( .A1(\mreg/_01142_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04648_ ), .ZN(\mreg/_01663_ ) );
INV_X1 \mreg/_07545_ ( .A(\mreg/_00041_ ), .ZN(\mreg/_01664_ ) );
AOI21_X1 \mreg/_07546_ ( .A(\mreg/_01663_ ), .B1(\mreg/_01664_ ), .B2(\mreg/_01173_ ), .ZN(\mreg/_01665_ ) );
AND4_X1 \mreg/_07547_ ( .A1(\mreg/_01656_ ), .A2(\mreg/_01661_ ), .A3(\mreg/_01662_ ), .A4(\mreg/_01665_ ), .ZN(\mreg/_01666_ ) );
BUF_X4 \mreg/_07548_ ( .A(\mreg/_01188_ ), .Z(\mreg/_01667_ ) );
NAND4_X1 \mreg/_07549_ ( .A1(\mreg/_01667_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04200_ ), .A4(\mreg/_01212_ ), .ZN(\mreg/_01668_ ) );
INV_X1 \mreg/_07550_ ( .A(\mreg/_04232_ ), .ZN(\mreg/_01669_ ) );
OAI21_X1 \mreg/_07551_ ( .A(\mreg/_01668_ ), .B1(\mreg/_01069_ ), .B2(\mreg/_01669_ ), .ZN(\mreg/_01670_ ) );
AOI221_X4 \mreg/_07552_ ( .A(\mreg/_01670_ ), .B1(\mreg/_04168_ ), .B2(\mreg/_01075_ ), .C1(\mreg/_04136_ ), .C2(\mreg/_01080_ ), .ZN(\mreg/_01671_ ) );
NAND3_X1 \mreg/_07553_ ( .A1(\mreg/_01091_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04360_ ), .ZN(\mreg/_01672_ ) );
NAND3_X1 \mreg/_07554_ ( .A1(\mreg/_01380_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04392_ ), .ZN(\mreg/_01673_ ) );
NAND2_X1 \mreg/_07555_ ( .A1(\mreg/_01672_ ), .A2(\mreg/_01673_ ), .ZN(\mreg/_01674_ ) );
AOI221_X4 \mreg/_07556_ ( .A(\mreg/_01674_ ), .B1(\mreg/_04328_ ), .B2(\mreg/_01205_ ), .C1(\mreg/_04296_ ), .C2(\mreg/_01207_ ), .ZN(\mreg/_01675_ ) );
NAND4_X1 \mreg/_07557_ ( .A1(\mreg/_01655_ ), .A2(\mreg/_01666_ ), .A3(\mreg/_01671_ ), .A4(\mreg/_01675_ ), .ZN(\mreg/_03912_ ) );
NAND3_X1 \mreg/_07558_ ( .A1(\mreg/_01084_ ), .A2(\mreg/_04553_ ), .A3(\mreg/_01299_ ), .ZN(\mreg/_01676_ ) );
NAND4_X1 \mreg/_07559_ ( .A1(\mreg/_01318_ ), .A2(\mreg/_01453_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04489_ ), .ZN(\mreg/_01677_ ) );
BUF_X4 \mreg/_07560_ ( .A(\mreg/_01190_ ), .Z(\mreg/_01678_ ) );
INV_X1 \mreg/_07561_ ( .A(\mreg/_04521_ ), .ZN(\mreg/_01679_ ) );
OAI21_X1 \mreg/_07562_ ( .A(\mreg/_01677_ ), .B1(\mreg/_01678_ ), .B2(\mreg/_01679_ ), .ZN(\mreg/_01680_ ) );
AOI221_X4 \mreg/_07563_ ( .A(\mreg/_01680_ ), .B1(\mreg/_04457_ ), .B2(\mreg/_01412_ ), .C1(\mreg/_04425_ ), .C2(\mreg/_01198_ ), .ZN(\mreg/_01681_ ) );
NAND3_X1 \mreg/_07564_ ( .A1(\mreg/_01305_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04585_ ), .ZN(\mreg/_01682_ ) );
AND3_X1 \mreg/_07565_ ( .A1(\mreg/_01143_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04649_ ), .ZN(\mreg/_01683_ ) );
INV_X1 \mreg/_07566_ ( .A(\mreg/_00042_ ), .ZN(\mreg/_01684_ ) );
AOI21_X1 \mreg/_07567_ ( .A(\mreg/_01683_ ), .B1(\mreg/_01684_ ), .B2(\mreg/_01173_ ), .ZN(\mreg/_01685_ ) );
AND4_X4 \mreg/_07568_ ( .A1(\mreg/_01676_ ), .A2(\mreg/_01681_ ), .A3(\mreg/_01682_ ), .A4(\mreg/_01685_ ), .ZN(\mreg/_01686_ ) );
NAND4_X1 \mreg/_07569_ ( .A1(\mreg/_01667_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04201_ ), .A4(\mreg/_01212_ ), .ZN(\mreg/_01687_ ) );
INV_X1 \mreg/_07570_ ( .A(\mreg/_04233_ ), .ZN(\mreg/_01688_ ) );
OAI21_X1 \mreg/_07571_ ( .A(\mreg/_01687_ ), .B1(\mreg/_01069_ ), .B2(\mreg/_01688_ ), .ZN(\mreg/_01689_ ) );
AOI221_X4 \mreg/_07572_ ( .A(\mreg/_01689_ ), .B1(\mreg/_04169_ ), .B2(\mreg/_01075_ ), .C1(\mreg/_04137_ ), .C2(\mreg/_01080_ ), .ZN(\mreg/_01690_ ) );
NAND3_X1 \mreg/_07573_ ( .A1(\mreg/_01092_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04361_ ), .ZN(\mreg/_01691_ ) );
NAND3_X1 \mreg/_07574_ ( .A1(\mreg/_01380_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04393_ ), .ZN(\mreg/_01692_ ) );
NAND2_X1 \mreg/_07575_ ( .A1(\mreg/_01691_ ), .A2(\mreg/_01692_ ), .ZN(\mreg/_01693_ ) );
AOI221_X4 \mreg/_07576_ ( .A(\mreg/_01693_ ), .B1(\mreg/_04329_ ), .B2(\mreg/_01205_ ), .C1(\mreg/_04297_ ), .C2(\mreg/_01207_ ), .ZN(\mreg/_01694_ ) );
AND3_X1 \mreg/_07577_ ( .A1(\mreg/_01072_ ), .A2(\mreg/_01103_ ), .A3(\mreg/_04265_ ), .ZN(\mreg/_01695_ ) );
AOI221_X4 \mreg/_07578_ ( .A(\mreg/_01695_ ), .B1(\mreg/_01106_ ), .B2(\mreg/_04713_ ), .C1(\mreg/_04617_ ), .C2(\mreg/_01221_ ), .ZN(\mreg/_01696_ ) );
AND3_X1 \mreg/_07579_ ( .A1(\mreg/_01092_ ), .A2(\mreg/_01144_ ), .A3(\mreg/_04809_ ), .ZN(\mreg/_01697_ ) );
AND3_X1 \mreg/_07580_ ( .A1(\mreg/_01097_ ), .A2(\mreg/_01122_ ), .A3(\mreg/_04841_ ), .ZN(\mreg/_01698_ ) );
AND3_X1 \mreg/_07581_ ( .A1(\mreg/_01058_ ), .A2(\mreg/_01122_ ), .A3(\mreg/_04777_ ), .ZN(\mreg/_01699_ ) );
AND3_X1 \mreg/_07582_ ( .A1(\mreg/_01126_ ), .A2(\mreg/_04745_ ), .A3(\mreg/_01086_ ), .ZN(\mreg/_01700_ ) );
NOR4_X1 \mreg/_07583_ ( .A1(\mreg/_01697_ ), .A2(\mreg/_01698_ ), .A3(\mreg/_01699_ ), .A4(\mreg/_01700_ ), .ZN(\mreg/_01701_ ) );
AND3_X1 \mreg/_07584_ ( .A1(\mreg/_01112_ ), .A2(\mreg/_01133_ ), .A3(\mreg/_03977_ ), .ZN(\mreg/_01702_ ) );
AND3_X1 \mreg/_07585_ ( .A1(\mreg/_01117_ ), .A2(\mreg/_01122_ ), .A3(\mreg/_03945_ ), .ZN(\mreg/_01703_ ) );
AND3_X1 \mreg/_07586_ ( .A1(\mreg/_01121_ ), .A2(\mreg/_01122_ ), .A3(\mreg/_04905_ ), .ZN(\mreg/_01704_ ) );
AND3_X1 \mreg/_07587_ ( .A1(\mreg/_01125_ ), .A2(\mreg/_04873_ ), .A3(\mreg/_01127_ ), .ZN(\mreg/_01705_ ) );
NOR4_X1 \mreg/_07588_ ( .A1(\mreg/_01702_ ), .A2(\mreg/_01703_ ), .A3(\mreg/_01704_ ), .A4(\mreg/_01705_ ), .ZN(\mreg/_01706_ ) );
NAND3_X1 \mreg/_07589_ ( .A1(\mreg/_01338_ ), .A2(\mreg/_04009_ ), .A3(\mreg/_01151_ ), .ZN(\mreg/_01707_ ) );
NAND3_X1 \mreg/_07590_ ( .A1(\mreg/_01142_ ), .A2(\mreg/_01217_ ), .A3(\mreg/_04073_ ), .ZN(\mreg/_01708_ ) );
NAND3_X1 \mreg/_07591_ ( .A1(\mreg/_01148_ ), .A2(\mreg/_01217_ ), .A3(\mreg/_04041_ ), .ZN(\mreg/_01709_ ) );
NAND3_X1 \mreg/_07592_ ( .A1(\mreg/_01140_ ), .A2(\mreg/_01118_ ), .A3(\mreg/_04105_ ), .ZN(\mreg/_01710_ ) );
AND4_X1 \mreg/_07593_ ( .A1(\mreg/_01707_ ), .A2(\mreg/_01708_ ), .A3(\mreg/_01709_ ), .A4(\mreg/_01710_ ), .ZN(\mreg/_01711_ ) );
AND4_X1 \mreg/_07594_ ( .A1(\mreg/_01696_ ), .A2(\mreg/_01701_ ), .A3(\mreg/_01706_ ), .A4(\mreg/_01711_ ), .ZN(\mreg/_01712_ ) );
NAND4_X1 \mreg/_07595_ ( .A1(\mreg/_01686_ ), .A2(\mreg/_01690_ ), .A3(\mreg/_01694_ ), .A4(\mreg/_01712_ ), .ZN(\mreg/_03913_ ) );
NAND3_X1 \mreg/_07596_ ( .A1(\mreg/_01083_ ), .A2(\mreg/_04554_ ), .A3(\mreg/_01597_ ), .ZN(\mreg/_01713_ ) );
NAND3_X1 \mreg/_07597_ ( .A1(\mreg/_01180_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04650_ ), .ZN(\mreg/_01714_ ) );
NAND3_X1 \mreg/_07598_ ( .A1(\mreg/_01182_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04586_ ), .ZN(\mreg/_01715_ ) );
INV_X1 \mreg/_07599_ ( .A(\mreg/_00043_ ), .ZN(\mreg/_01716_ ) );
NAND3_X1 \mreg/_07600_ ( .A1(\mreg/_01184_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_01716_ ), .ZN(\mreg/_01717_ ) );
AND4_X1 \mreg/_07601_ ( .A1(\mreg/_01713_ ), .A2(\mreg/_01714_ ), .A3(\mreg/_01715_ ), .A4(\mreg/_01717_ ), .ZN(\mreg/_01718_ ) );
AND3_X1 \mreg/_07602_ ( .A1(\mreg/_01077_ ), .A2(\mreg/_04426_ ), .A3(\mreg/_01127_ ), .ZN(\mreg/_01719_ ) );
NAND4_X1 \mreg/_07603_ ( .A1(\mreg/_01188_ ), .A2(\mreg/_01161_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04490_ ), .ZN(\mreg/_01720_ ) );
INV_X1 \mreg/_07604_ ( .A(\mreg/_04522_ ), .ZN(\mreg/_01721_ ) );
OAI21_X1 \mreg/_07605_ ( .A(\mreg/_01720_ ), .B1(\mreg/_01191_ ), .B2(\mreg/_01721_ ), .ZN(\mreg/_01722_ ) );
AOI211_X4 \mreg/_07606_ ( .A(\mreg/_01719_ ), .B(\mreg/_01722_ ), .C1(\mreg/_04458_ ), .C2(\mreg/_01196_ ), .ZN(\mreg/_01723_ ) );
NAND3_X1 \mreg/_07607_ ( .A1(\mreg/_01323_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04362_ ), .ZN(\mreg/_01724_ ) );
NAND3_X1 \mreg/_07608_ ( .A1(\mreg/_01496_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04394_ ), .ZN(\mreg/_01725_ ) );
NAND2_X1 \mreg/_07609_ ( .A1(\mreg/_01724_ ), .A2(\mreg/_01725_ ), .ZN(\mreg/_01726_ ) );
AOI221_X4 \mreg/_07610_ ( .A(\mreg/_01726_ ), .B1(\mreg/_04330_ ), .B2(\mreg/_01611_ ), .C1(\mreg/_04298_ ), .C2(\mreg/_01499_ ), .ZN(\mreg/_01727_ ) );
NAND4_X1 \mreg/_07611_ ( .A1(\mreg/_01501_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04202_ ), .A4(\mreg/_01372_ ), .ZN(\mreg/_01728_ ) );
INV_X1 \mreg/_07612_ ( .A(\mreg/_04234_ ), .ZN(\mreg/_01729_ ) );
OAI21_X1 \mreg/_07613_ ( .A(\mreg/_01728_ ), .B1(\mreg/_01374_ ), .B2(\mreg/_01729_ ), .ZN(\mreg/_01730_ ) );
AOI221_X4 \mreg/_07614_ ( .A(\mreg/_01730_ ), .B1(\mreg/_04170_ ), .B2(\mreg/_01465_ ), .C1(\mreg/_04138_ ), .C2(\mreg/_01505_ ), .ZN(\mreg/_01731_ ) );
AND4_X4 \mreg/_07615_ ( .A1(\mreg/_01718_ ), .A2(\mreg/_01723_ ), .A3(\mreg/_01727_ ), .A4(\mreg/_01731_ ), .ZN(\mreg/_01732_ ) );
NAND3_X1 \mreg/_07616_ ( .A1(\mreg/_01275_ ), .A2(\mreg/_01277_ ), .A3(\mreg/_04810_ ), .ZN(\mreg/_01733_ ) );
AND3_X1 \mreg/_07617_ ( .A1(\mreg/_01072_ ), .A2(\mreg/_01103_ ), .A3(\mreg/_04266_ ), .ZN(\mreg/_01734_ ) );
AOI221_X4 \mreg/_07618_ ( .A(\mreg/_01734_ ), .B1(\mreg/_01106_ ), .B2(\mreg/_04714_ ), .C1(\mreg/_04618_ ), .C2(\mreg/_01221_ ), .ZN(\mreg/_01735_ ) );
NAND3_X1 \mreg/_07619_ ( .A1(\mreg/_01281_ ), .A2(\mreg/_01282_ ), .A3(\mreg/_04842_ ), .ZN(\mreg/_01736_ ) );
AOI22_X1 \mreg/_07620_ ( .A1(\mreg/_01284_ ), .A2(\mreg/_04778_ ), .B1(\mreg/_04746_ ), .B2(\mreg/_01230_ ), .ZN(\mreg/_01737_ ) );
AND4_X1 \mreg/_07621_ ( .A1(\mreg/_01733_ ), .A2(\mreg/_01735_ ), .A3(\mreg/_01736_ ), .A4(\mreg/_01737_ ), .ZN(\mreg/_01738_ ) );
NAND3_X1 \mreg/_07622_ ( .A1(\mreg/_01156_ ), .A2(\mreg/_01287_ ), .A3(\mreg/_04906_ ), .ZN(\mreg/_01739_ ) );
NAND3_X1 \mreg/_07623_ ( .A1(\mreg/_01159_ ), .A2(\mreg/_01289_ ), .A3(\mreg/_03946_ ), .ZN(\mreg/_01740_ ) );
NAND3_X1 \mreg/_07624_ ( .A1(\mreg/_01292_ ), .A2(\mreg/_01293_ ), .A3(\mreg/_04874_ ), .ZN(\mreg/_01741_ ) );
NAND3_X1 \mreg/_07625_ ( .A1(\mreg/_01165_ ), .A2(\mreg/_01477_ ), .A3(\mreg/_03978_ ), .ZN(\mreg/_01742_ ) );
AND4_X1 \mreg/_07626_ ( .A1(\mreg/_01739_ ), .A2(\mreg/_01740_ ), .A3(\mreg/_01741_ ), .A4(\mreg/_01742_ ), .ZN(\mreg/_01743_ ) );
NAND3_X1 \mreg/_07627_ ( .A1(\mreg/_01298_ ), .A2(\mreg/_04010_ ), .A3(\mreg/_01299_ ), .ZN(\mreg/_01744_ ) );
NAND3_X1 \mreg/_07628_ ( .A1(\mreg/_01301_ ), .A2(\mreg/_01302_ ), .A3(\mreg/_04074_ ), .ZN(\mreg/_01745_ ) );
NAND3_X1 \mreg/_07629_ ( .A1(\mreg/_01305_ ), .A2(\mreg/_01295_ ), .A3(\mreg/_04042_ ), .ZN(\mreg/_01746_ ) );
NAND3_X1 \mreg/_07630_ ( .A1(\mreg/_01308_ ), .A2(\mreg/_01309_ ), .A3(\mreg/_04106_ ), .ZN(\mreg/_01747_ ) );
AND4_X1 \mreg/_07631_ ( .A1(\mreg/_01744_ ), .A2(\mreg/_01745_ ), .A3(\mreg/_01746_ ), .A4(\mreg/_01747_ ), .ZN(\mreg/_01748_ ) );
NAND4_X1 \mreg/_07632_ ( .A1(\mreg/_01732_ ), .A2(\mreg/_01738_ ), .A3(\mreg/_01743_ ), .A4(\mreg/_01748_ ), .ZN(\mreg/_03914_ ) );
NAND3_X1 \mreg/_07633_ ( .A1(\mreg/_01147_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04587_ ), .ZN(\mreg/_01749_ ) );
NAND3_X1 \mreg/_07634_ ( .A1(\mreg/_01255_ ), .A2(\mreg/_04555_ ), .A3(\mreg/_01150_ ), .ZN(\mreg/_01750_ ) );
NAND2_X1 \mreg/_07635_ ( .A1(\mreg/_01749_ ), .A2(\mreg/_01750_ ), .ZN(\mreg/_01751_ ) );
INV_X1 \mreg/_07636_ ( .A(\mreg/_00044_ ), .ZN(\mreg/_01752_ ) );
AOI221_X1 \mreg/_07637_ ( .A(\mreg/_01751_ ), .B1(\mreg/_01752_ ), .B2(\mreg/_01173_ ), .C1(\mreg/_04651_ ), .C2(\mreg/_01175_ ), .ZN(\mreg/_01753_ ) );
NAND4_X1 \mreg/_07638_ ( .A1(\mreg/_01318_ ), .A2(\mreg/_01453_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04491_ ), .ZN(\mreg/_01754_ ) );
INV_X1 \mreg/_07639_ ( .A(\mreg/_04523_ ), .ZN(\mreg/_01755_ ) );
OAI21_X1 \mreg/_07640_ ( .A(\mreg/_01754_ ), .B1(\mreg/_01678_ ), .B2(\mreg/_01755_ ), .ZN(\mreg/_01756_ ) );
AOI221_X4 \mreg/_07641_ ( .A(\mreg/_01756_ ), .B1(\mreg/_04459_ ), .B2(\mreg/_01412_ ), .C1(\mreg/_04427_ ), .C2(\mreg/_01198_ ), .ZN(\mreg/_01757_ ) );
NAND3_X1 \mreg/_07642_ ( .A1(\mreg/_01323_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04363_ ), .ZN(\mreg/_01758_ ) );
NAND3_X1 \mreg/_07643_ ( .A1(\mreg/_01496_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04395_ ), .ZN(\mreg/_01759_ ) );
NAND2_X1 \mreg/_07644_ ( .A1(\mreg/_01758_ ), .A2(\mreg/_01759_ ), .ZN(\mreg/_01760_ ) );
AOI221_X4 \mreg/_07645_ ( .A(\mreg/_01760_ ), .B1(\mreg/_04331_ ), .B2(\mreg/_01611_ ), .C1(\mreg/_04299_ ), .C2(\mreg/_01499_ ), .ZN(\mreg/_01761_ ) );
NAND4_X1 \mreg/_07646_ ( .A1(\mreg/_01188_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04203_ ), .A4(\mreg/_01209_ ), .ZN(\mreg/_01762_ ) );
NAND4_X1 \mreg/_07647_ ( .A1(\mreg/_01211_ ), .A2(\mreg/_01212_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04235_ ), .ZN(\mreg/_01763_ ) );
NAND2_X1 \mreg/_07648_ ( .A1(\mreg/_01762_ ), .A2(\mreg/_01763_ ), .ZN(\mreg/_01764_ ) );
AOI221_X4 \mreg/_07649_ ( .A(\mreg/_01764_ ), .B1(\mreg/_01079_ ), .B2(\mreg/_04139_ ), .C1(\mreg/_04171_ ), .C2(\mreg/_01075_ ), .ZN(\mreg/_01765_ ) );
AND4_X4 \mreg/_07650_ ( .A1(\mreg/_01753_ ), .A2(\mreg/_01757_ ), .A3(\mreg/_01761_ ), .A4(\mreg/_01765_ ), .ZN(\mreg/_01766_ ) );
AND3_X1 \mreg/_07651_ ( .A1(\mreg/_01107_ ), .A2(\mreg/_01217_ ), .A3(\mreg/_04267_ ), .ZN(\mreg/_01767_ ) );
AOI221_X4 \mreg/_07652_ ( .A(\mreg/_01767_ ), .B1(\mreg/_01219_ ), .B2(\mreg/_04715_ ), .C1(\mreg/_04619_ ), .C2(\mreg/_01222_ ), .ZN(\mreg/_01768_ ) );
NAND3_X1 \mreg/_07653_ ( .A1(\mreg/_01059_ ), .A2(\mreg/_01287_ ), .A3(\mreg/_04779_ ), .ZN(\mreg/_01769_ ) );
NAND3_X1 \mreg/_07654_ ( .A1(\mreg/_01275_ ), .A2(\mreg/_01289_ ), .A3(\mreg/_04811_ ), .ZN(\mreg/_01770_ ) );
NAND3_X1 \mreg/_07655_ ( .A1(\mreg/_01281_ ), .A2(\mreg/_01306_ ), .A3(\mreg/_04843_ ), .ZN(\mreg/_01771_ ) );
NAND3_X1 \mreg/_07656_ ( .A1(\mreg/_01339_ ), .A2(\mreg/_01087_ ), .A3(\mreg/_04747_ ), .ZN(\mreg/_01772_ ) );
AND4_X1 \mreg/_07657_ ( .A1(\mreg/_01769_ ), .A2(\mreg/_01770_ ), .A3(\mreg/_01771_ ), .A4(\mreg/_01772_ ), .ZN(\mreg/_01773_ ) );
NAND3_X1 \mreg/_07658_ ( .A1(\mreg/_01301_ ), .A2(\mreg/_01289_ ), .A3(\mreg/_04075_ ), .ZN(\mreg/_01774_ ) );
NAND3_X1 \mreg/_07659_ ( .A1(\mreg/_01121_ ), .A2(\mreg/_01130_ ), .A3(\mreg/_04907_ ), .ZN(\mreg/_01775_ ) );
NAND3_X1 \mreg/_07660_ ( .A1(\mreg/_01158_ ), .A2(\mreg/_01144_ ), .A3(\mreg/_03947_ ), .ZN(\mreg/_01776_ ) );
NAND3_X1 \mreg/_07661_ ( .A1(\mreg/_01338_ ), .A2(\mreg/_01162_ ), .A3(\mreg/_04875_ ), .ZN(\mreg/_01777_ ) );
NAND3_X1 \mreg/_07662_ ( .A1(\mreg/_01112_ ), .A2(\mreg/_01217_ ), .A3(\mreg/_03979_ ), .ZN(\mreg/_01778_ ) );
AND4_X1 \mreg/_07663_ ( .A1(\mreg/_01775_ ), .A2(\mreg/_01776_ ), .A3(\mreg/_01777_ ), .A4(\mreg/_01778_ ), .ZN(\mreg/_01779_ ) );
NAND3_X1 \mreg/_07664_ ( .A1(\mreg/_01308_ ), .A2(\mreg/_01295_ ), .A3(\mreg/_04107_ ), .ZN(\mreg/_01780_ ) );
AND3_X1 \mreg/_07665_ ( .A1(\mreg/_01148_ ), .A2(\mreg/_01622_ ), .A3(\mreg/_04043_ ), .ZN(\mreg/_01781_ ) );
AND3_X1 \mreg/_07666_ ( .A1(\mreg/_01338_ ), .A2(\mreg/_04011_ ), .A3(\mreg/_01151_ ), .ZN(\mreg/_01782_ ) );
NOR2_X1 \mreg/_07667_ ( .A1(\mreg/_01781_ ), .A2(\mreg/_01782_ ), .ZN(\mreg/_01783_ ) );
AND4_X1 \mreg/_07668_ ( .A1(\mreg/_01774_ ), .A2(\mreg/_01779_ ), .A3(\mreg/_01780_ ), .A4(\mreg/_01783_ ), .ZN(\mreg/_01784_ ) );
NAND4_X1 \mreg/_07669_ ( .A1(\mreg/_01766_ ), .A2(\mreg/_01768_ ), .A3(\mreg/_01773_ ), .A4(\mreg/_01784_ ), .ZN(\mreg/_03915_ ) );
NAND3_X1 \mreg/_07670_ ( .A1(\mreg/_01125_ ), .A2(\mreg/_01086_ ), .A3(\mreg/_04748_ ), .ZN(\mreg/_01785_ ) );
INV_X4 \mreg/_07671_ ( .A(\mreg/_01105_ ), .ZN(\mreg/_01786_ ) );
INV_X1 \mreg/_07672_ ( .A(\mreg/_04716_ ), .ZN(\mreg/_01787_ ) );
OAI21_X1 \mreg/_07673_ ( .A(\mreg/_01785_ ), .B1(\mreg/_01786_ ), .B2(\mreg/_01787_ ), .ZN(\mreg/_01788_ ) );
AOI221_X4 \mreg/_07674_ ( .A(\mreg/_01788_ ), .B1(\mreg/_04812_ ), .B2(\mreg/_01430_ ), .C1(\mreg/_04780_ ), .C2(\mreg/_01228_ ), .ZN(\mreg/_01789_ ) );
NAND3_X1 \mreg/_07675_ ( .A1(\mreg/_01139_ ), .A2(\mreg/_01357_ ), .A3(\mreg/_04108_ ), .ZN(\mreg/_01790_ ) );
NAND2_X1 \mreg/_07676_ ( .A1(\mreg/_01146_ ), .A2(\mreg/_01108_ ), .ZN(\mreg/_01791_ ) );
INV_X1 \mreg/_07677_ ( .A(\mreg/_04044_ ), .ZN(\mreg/_01792_ ) );
OAI21_X1 \mreg/_07678_ ( .A(\mreg/_01790_ ), .B1(\mreg/_01791_ ), .B2(\mreg/_01792_ ), .ZN(\mreg/_01793_ ) );
AOI221_X4 \mreg/_07679_ ( .A(\mreg/_01793_ ), .B1(\mreg/_03948_ ), .B2(\mreg/_01361_ ), .C1(\mreg/_04908_ ), .C2(\mreg/_01363_ ), .ZN(\mreg/_01794_ ) );
NAND4_X1 \mreg/_07680_ ( .A1(\mreg/_01269_ ), .A2(\mreg/_01366_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04492_ ), .ZN(\mreg/_01795_ ) );
INV_X1 \mreg/_07681_ ( .A(\mreg/_04524_ ), .ZN(\mreg/_01796_ ) );
OAI21_X1 \mreg/_07682_ ( .A(\mreg/_01795_ ), .B1(\mreg/_01190_ ), .B2(\mreg/_01796_ ), .ZN(\mreg/_01797_ ) );
INV_X1 \mreg/_07683_ ( .A(\mreg/_00045_ ), .ZN(\mreg/_01798_ ) );
AOI221_X4 \mreg/_07684_ ( .A(\mreg/_01797_ ), .B1(\mreg/_01798_ ), .B2(\mreg/_01172_ ), .C1(\mreg/_04652_ ), .C2(\mreg/_01175_ ), .ZN(\mreg/_01799_ ) );
NAND4_X1 \mreg/_07685_ ( .A1(\mreg/_01501_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04204_ ), .A4(\mreg/_01372_ ), .ZN(\mreg/_01800_ ) );
INV_X1 \mreg/_07686_ ( .A(\mreg/_04236_ ), .ZN(\mreg/_01801_ ) );
OAI21_X1 \mreg/_07687_ ( .A(\mreg/_01800_ ), .B1(\mreg/_01374_ ), .B2(\mreg/_01801_ ), .ZN(\mreg/_01802_ ) );
AOI221_X4 \mreg/_07688_ ( .A(\mreg/_01802_ ), .B1(\mreg/_04332_ ), .B2(\mreg/_01204_ ), .C1(\mreg/_04300_ ), .C2(\mreg/_01377_ ), .ZN(\mreg/_01803_ ) );
AND4_X4 \mreg/_07689_ ( .A1(\mreg/_01789_ ), .A2(\mreg/_01794_ ), .A3(\mreg/_01799_ ), .A4(\mreg/_01803_ ), .ZN(\mreg/_01804_ ) );
NAND3_X1 \mreg/_07690_ ( .A1(\mreg/_01339_ ), .A2(\mreg/_04012_ ), .A3(\mreg/_01242_ ), .ZN(\mreg/_01805_ ) );
INV_X1 \mreg/_07691_ ( .A(\mreg/_04076_ ), .ZN(\mreg/_01806_ ) );
INV_X1 \mreg/_07692_ ( .A(\mreg/_03980_ ), .ZN(\mreg/_01807_ ) );
OAI221_X1 \mreg/_07693_ ( .A(\mreg/_01805_ ), .B1(\mreg/_01393_ ), .B2(\mreg/_01806_ ), .C1(\mreg/_01807_ ), .C2(\mreg/_01396_ ), .ZN(\mreg/_01808_ ) );
AND3_X1 \mreg/_07694_ ( .A1(\mreg/_01381_ ), .A2(\mreg/_01233_ ), .A3(\mreg/_04844_ ), .ZN(\mreg/_01809_ ) );
AND3_X1 \mreg/_07695_ ( .A1(\mreg/_01241_ ), .A2(\mreg/_04876_ ), .A3(\mreg/_01163_ ), .ZN(\mreg/_01810_ ) );
NAND3_X1 \mreg/_07696_ ( .A1(\mreg/_01383_ ), .A2(\mreg/_01384_ ), .A3(\mreg/_04268_ ), .ZN(\mreg/_01811_ ) );
NAND3_X1 \mreg/_07697_ ( .A1(\mreg/_01386_ ), .A2(\mreg/_01387_ ), .A3(\mreg/_04620_ ), .ZN(\mreg/_01812_ ) );
NAND2_X1 \mreg/_07698_ ( .A1(\mreg/_01811_ ), .A2(\mreg/_01812_ ), .ZN(\mreg/_01813_ ) );
NOR4_X1 \mreg/_07699_ ( .A1(\mreg/_01808_ ), .A2(\mreg/_01809_ ), .A3(\mreg/_01810_ ), .A4(\mreg/_01813_ ), .ZN(\mreg/_01814_ ) );
NAND3_X1 \mreg/_07700_ ( .A1(\mreg/_01156_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04460_ ), .ZN(\mreg/_01815_ ) );
NAND3_X1 \mreg/_07701_ ( .A1(\mreg/_01305_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04588_ ), .ZN(\mreg/_01816_ ) );
NAND3_X1 \mreg/_07702_ ( .A1(\mreg/_01084_ ), .A2(\mreg/_04556_ ), .A3(\mreg/_01242_ ), .ZN(\mreg/_01817_ ) );
NAND3_X1 \mreg/_07703_ ( .A1(\mreg/_01084_ ), .A2(\mreg/_04428_ ), .A3(\mreg/_01163_ ), .ZN(\mreg/_01818_ ) );
AND4_X1 \mreg/_07704_ ( .A1(\mreg/_01815_ ), .A2(\mreg/_01816_ ), .A3(\mreg/_01817_ ), .A4(\mreg/_01818_ ), .ZN(\mreg/_01819_ ) );
NAND3_X1 \mreg/_07705_ ( .A1(\mreg/_01091_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04364_ ), .ZN(\mreg/_01820_ ) );
NAND3_X1 \mreg/_07706_ ( .A1(\mreg/_01380_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04396_ ), .ZN(\mreg/_01821_ ) );
NAND2_X1 \mreg/_07707_ ( .A1(\mreg/_01820_ ), .A2(\mreg/_01821_ ), .ZN(\mreg/_01822_ ) );
AOI221_X4 \mreg/_07708_ ( .A(\mreg/_01822_ ), .B1(\mreg/_04172_ ), .B2(\mreg/_01075_ ), .C1(\mreg/_04140_ ), .C2(\mreg/_01080_ ), .ZN(\mreg/_01823_ ) );
NAND4_X1 \mreg/_07709_ ( .A1(\mreg/_01804_ ), .A2(\mreg/_01814_ ), .A3(\mreg/_01819_ ), .A4(\mreg/_01823_ ), .ZN(\mreg/_03916_ ) );
NAND3_X1 \mreg/_07710_ ( .A1(\mreg/_01125_ ), .A2(\mreg/_01086_ ), .A3(\mreg/_04749_ ), .ZN(\mreg/_01824_ ) );
INV_X1 \mreg/_07711_ ( .A(\mreg/_04717_ ), .ZN(\mreg/_01825_ ) );
OAI21_X1 \mreg/_07712_ ( .A(\mreg/_01824_ ), .B1(\mreg/_01786_ ), .B2(\mreg/_01825_ ), .ZN(\mreg/_01826_ ) );
AOI221_X4 \mreg/_07713_ ( .A(\mreg/_01826_ ), .B1(\mreg/_04813_ ), .B2(\mreg/_01430_ ), .C1(\mreg/_04781_ ), .C2(\mreg/_01228_ ), .ZN(\mreg/_01827_ ) );
NAND3_X1 \mreg/_07714_ ( .A1(\mreg/_01139_ ), .A2(\mreg/_01108_ ), .A3(\mreg/_04109_ ), .ZN(\mreg/_01828_ ) );
INV_X1 \mreg/_07715_ ( .A(\mreg/_04045_ ), .ZN(\mreg/_01829_ ) );
OAI21_X1 \mreg/_07716_ ( .A(\mreg/_01828_ ), .B1(\mreg/_01791_ ), .B2(\mreg/_01829_ ), .ZN(\mreg/_01830_ ) );
AOI221_X1 \mreg/_07717_ ( .A(\mreg/_01830_ ), .B1(\mreg/_03949_ ), .B2(\mreg/_01361_ ), .C1(\mreg/_04909_ ), .C2(\mreg/_01363_ ), .ZN(\mreg/_01831_ ) );
NAND4_X1 \mreg/_07718_ ( .A1(\mreg/_01365_ ), .A2(\mreg/_01366_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04493_ ), .ZN(\mreg/_01832_ ) );
INV_X1 \mreg/_07719_ ( .A(\mreg/_04525_ ), .ZN(\mreg/_01833_ ) );
OAI21_X1 \mreg/_07720_ ( .A(\mreg/_01832_ ), .B1(\mreg/_01190_ ), .B2(\mreg/_01833_ ), .ZN(\mreg/_01834_ ) );
INV_X1 \mreg/_07721_ ( .A(\mreg/_00046_ ), .ZN(\mreg/_01835_ ) );
AOI221_X1 \mreg/_07722_ ( .A(\mreg/_01834_ ), .B1(\mreg/_01835_ ), .B2(\mreg/_01172_ ), .C1(\mreg/_04653_ ), .C2(\mreg/_01174_ ), .ZN(\mreg/_01836_ ) );
NAND4_X1 \mreg/_07723_ ( .A1(\mreg/_01089_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04205_ ), .A4(\mreg/_01062_ ), .ZN(\mreg/_01837_ ) );
INV_X1 \mreg/_07724_ ( .A(\mreg/_04237_ ), .ZN(\mreg/_01838_ ) );
OAI21_X1 \mreg/_07725_ ( .A(\mreg/_01837_ ), .B1(\mreg/_01068_ ), .B2(\mreg/_01838_ ), .ZN(\mreg/_01839_ ) );
AOI221_X4 \mreg/_07726_ ( .A(\mreg/_01839_ ), .B1(\mreg/_04333_ ), .B2(\mreg/_01204_ ), .C1(\mreg/_04301_ ), .C2(\mreg/_01377_ ), .ZN(\mreg/_01840_ ) );
NAND4_X1 \mreg/_07727_ ( .A1(\mreg/_01827_ ), .A2(\mreg/_01831_ ), .A3(\mreg/_01836_ ), .A4(\mreg/_01840_ ), .ZN(\mreg/_01841_ ) );
NAND3_X1 \mreg/_07728_ ( .A1(\mreg/_01381_ ), .A2(\mreg/_01239_ ), .A3(\mreg/_04845_ ), .ZN(\mreg/_01842_ ) );
NAND3_X1 \mreg/_07729_ ( .A1(\mreg/_01383_ ), .A2(\mreg/_01384_ ), .A3(\mreg/_04269_ ), .ZN(\mreg/_01843_ ) );
NAND3_X1 \mreg/_07730_ ( .A1(\mreg/_01386_ ), .A2(\mreg/_01387_ ), .A3(\mreg/_04621_ ), .ZN(\mreg/_01844_ ) );
NAND3_X1 \mreg/_07731_ ( .A1(\mreg/_01241_ ), .A2(\mreg/_01163_ ), .A3(\mreg/_04877_ ), .ZN(\mreg/_01845_ ) );
NAND4_X1 \mreg/_07732_ ( .A1(\mreg/_01842_ ), .A2(\mreg/_01843_ ), .A3(\mreg/_01844_ ), .A4(\mreg/_01845_ ), .ZN(\mreg/_01846_ ) );
NAND3_X1 \mreg/_07733_ ( .A1(\mreg/_01291_ ), .A2(\mreg/_04013_ ), .A3(\mreg/_01391_ ), .ZN(\mreg/_01847_ ) );
INV_X1 \mreg/_07734_ ( .A(\mreg/_04077_ ), .ZN(\mreg/_01848_ ) );
INV_X1 \mreg/_07735_ ( .A(\mreg/_03981_ ), .ZN(\mreg/_01849_ ) );
OAI221_X1 \mreg/_07736_ ( .A(\mreg/_01847_ ), .B1(\mreg/_01393_ ), .B2(\mreg/_01848_ ), .C1(\mreg/_01849_ ), .C2(\mreg/_01396_ ), .ZN(\mreg/_01850_ ) );
NAND3_X2 \mreg/_07737_ ( .A1(\mreg/_01398_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04365_ ), .ZN(\mreg/_01851_ ) );
NAND3_X2 \mreg/_07738_ ( .A1(\mreg/_01096_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04397_ ), .ZN(\mreg/_01852_ ) );
NAND2_X1 \mreg/_07739_ ( .A1(\mreg/_01851_ ), .A2(\mreg/_01852_ ), .ZN(\mreg/_01853_ ) );
AOI221_X2 \mreg/_07740_ ( .A(\mreg/_01853_ ), .B1(\mreg/_04173_ ), .B2(\mreg/_01074_ ), .C1(\mreg/_04141_ ), .C2(\mreg/_01079_ ), .ZN(\mreg/_01854_ ) );
AND3_X1 \mreg/_07741_ ( .A1(\mreg/_01255_ ), .A2(\mreg/_04429_ ), .A3(\mreg/_01127_ ), .ZN(\mreg/_01855_ ) );
AOI21_X1 \mreg/_07742_ ( .A(\mreg/_01855_ ), .B1(\mreg/_01196_ ), .B2(\mreg/_04461_ ), .ZN(\mreg/_01856_ ) );
NAND3_X1 \mreg/_07743_ ( .A1(\mreg/_01177_ ), .A2(\mreg/_04557_ ), .A3(\mreg/_01178_ ), .ZN(\mreg/_01857_ ) );
NAND3_X1 \mreg/_07744_ ( .A1(\mreg/_01304_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04589_ ), .ZN(\mreg/_01858_ ) );
NAND4_X4 \mreg/_07745_ ( .A1(\mreg/_01854_ ), .A2(\mreg/_01856_ ), .A3(\mreg/_01857_ ), .A4(\mreg/_01858_ ), .ZN(\mreg/_01859_ ) );
OR4_X2 \mreg/_07746_ ( .A1(\mreg/_01841_ ), .A2(\mreg/_01846_ ), .A3(\mreg/_01850_ ), .A4(\mreg/_01859_ ), .ZN(\mreg/_03917_ ) );
NAND3_X1 \mreg/_07747_ ( .A1(\mreg/_01083_ ), .A2(\mreg/_04558_ ), .A3(\mreg/_01597_ ), .ZN(\mreg/_01860_ ) );
NAND3_X1 \mreg/_07748_ ( .A1(\mreg/_01180_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04654_ ), .ZN(\mreg/_01861_ ) );
NAND3_X1 \mreg/_07749_ ( .A1(\mreg/_01182_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04590_ ), .ZN(\mreg/_01862_ ) );
INV_X1 \mreg/_07750_ ( .A(\mreg/_00047_ ), .ZN(\mreg/_01863_ ) );
NAND3_X1 \mreg/_07751_ ( .A1(\mreg/_01184_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_01863_ ), .ZN(\mreg/_01864_ ) );
AND4_X1 \mreg/_07752_ ( .A1(\mreg/_01860_ ), .A2(\mreg/_01861_ ), .A3(\mreg/_01862_ ), .A4(\mreg/_01864_ ), .ZN(\mreg/_01865_ ) );
NAND4_X1 \mreg/_07753_ ( .A1(\mreg/_01318_ ), .A2(\mreg/_01453_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04494_ ), .ZN(\mreg/_01866_ ) );
INV_X1 \mreg/_07754_ ( .A(\mreg/_04526_ ), .ZN(\mreg/_01867_ ) );
OAI21_X1 \mreg/_07755_ ( .A(\mreg/_01866_ ), .B1(\mreg/_01678_ ), .B2(\mreg/_01867_ ), .ZN(\mreg/_01868_ ) );
AOI221_X4 \mreg/_07756_ ( .A(\mreg/_01868_ ), .B1(\mreg/_04462_ ), .B2(\mreg/_01412_ ), .C1(\mreg/_04430_ ), .C2(\mreg/_01198_ ), .ZN(\mreg/_01869_ ) );
NAND3_X1 \mreg/_07757_ ( .A1(\mreg/_01323_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04366_ ), .ZN(\mreg/_01870_ ) );
NAND3_X1 \mreg/_07758_ ( .A1(\mreg/_01496_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04398_ ), .ZN(\mreg/_01871_ ) );
NAND2_X1 \mreg/_07759_ ( .A1(\mreg/_01870_ ), .A2(\mreg/_01871_ ), .ZN(\mreg/_01872_ ) );
AOI221_X4 \mreg/_07760_ ( .A(\mreg/_01872_ ), .B1(\mreg/_04334_ ), .B2(\mreg/_01611_ ), .C1(\mreg/_04302_ ), .C2(\mreg/_01499_ ), .ZN(\mreg/_01873_ ) );
NAND4_X1 \mreg/_07761_ ( .A1(\mreg/_01501_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04206_ ), .A4(\mreg/_01372_ ), .ZN(\mreg/_01874_ ) );
INV_X1 \mreg/_07762_ ( .A(\mreg/_04238_ ), .ZN(\mreg/_01875_ ) );
OAI21_X1 \mreg/_07763_ ( .A(\mreg/_01874_ ), .B1(\mreg/_01374_ ), .B2(\mreg/_01875_ ), .ZN(\mreg/_01876_ ) );
AOI221_X4 \mreg/_07764_ ( .A(\mreg/_01876_ ), .B1(\mreg/_04174_ ), .B2(\mreg/_01465_ ), .C1(\mreg/_04142_ ), .C2(\mreg/_01505_ ), .ZN(\mreg/_01877_ ) );
AND4_X2 \mreg/_07765_ ( .A1(\mreg/_01865_ ), .A2(\mreg/_01869_ ), .A3(\mreg/_01873_ ), .A4(\mreg/_01877_ ), .ZN(\mreg/_01878_ ) );
NAND3_X1 \mreg/_07766_ ( .A1(\mreg/_01275_ ), .A2(\mreg/_01277_ ), .A3(\mreg/_04814_ ), .ZN(\mreg/_01879_ ) );
AND3_X1 \mreg/_07767_ ( .A1(\mreg/_01072_ ), .A2(\mreg/_01357_ ), .A3(\mreg/_04270_ ), .ZN(\mreg/_01880_ ) );
AOI221_X4 \mreg/_07768_ ( .A(\mreg/_01880_ ), .B1(\mreg/_01106_ ), .B2(\mreg/_04718_ ), .C1(\mreg/_04622_ ), .C2(\mreg/_01221_ ), .ZN(\mreg/_01881_ ) );
NAND3_X1 \mreg/_07769_ ( .A1(\mreg/_01281_ ), .A2(\mreg/_01302_ ), .A3(\mreg/_04846_ ), .ZN(\mreg/_01882_ ) );
AOI22_X1 \mreg/_07770_ ( .A1(\mreg/_01284_ ), .A2(\mreg/_04782_ ), .B1(\mreg/_04750_ ), .B2(\mreg/_01230_ ), .ZN(\mreg/_01883_ ) );
AND4_X1 \mreg/_07771_ ( .A1(\mreg/_01879_ ), .A2(\mreg/_01881_ ), .A3(\mreg/_01882_ ), .A4(\mreg/_01883_ ), .ZN(\mreg/_01884_ ) );
NAND3_X1 \mreg/_07772_ ( .A1(\mreg/_01156_ ), .A2(\mreg/_01436_ ), .A3(\mreg/_04910_ ), .ZN(\mreg/_01885_ ) );
NAND3_X1 \mreg/_07773_ ( .A1(\mreg/_01159_ ), .A2(\mreg/_01289_ ), .A3(\mreg/_03950_ ), .ZN(\mreg/_01886_ ) );
NAND3_X1 \mreg/_07774_ ( .A1(\mreg/_01292_ ), .A2(\mreg/_01293_ ), .A3(\mreg/_04878_ ), .ZN(\mreg/_01887_ ) );
NAND3_X1 \mreg/_07775_ ( .A1(\mreg/_01165_ ), .A2(\mreg/_01477_ ), .A3(\mreg/_03982_ ), .ZN(\mreg/_01888_ ) );
AND4_X1 \mreg/_07776_ ( .A1(\mreg/_01885_ ), .A2(\mreg/_01886_ ), .A3(\mreg/_01887_ ), .A4(\mreg/_01888_ ), .ZN(\mreg/_01889_ ) );
AND3_X1 \mreg/_07777_ ( .A1(\mreg/_01232_ ), .A2(\mreg/_01233_ ), .A3(\mreg/_04078_ ), .ZN(\mreg/_01890_ ) );
AND3_X1 \mreg/_07778_ ( .A1(\mreg/_01235_ ), .A2(\mreg/_01384_ ), .A3(\mreg/_04046_ ), .ZN(\mreg/_01891_ ) );
AND3_X1 \mreg/_07779_ ( .A1(\mreg/_01238_ ), .A2(\mreg/_01248_ ), .A3(\mreg/_04110_ ), .ZN(\mreg/_01892_ ) );
AND3_X1 \mreg/_07780_ ( .A1(\mreg/_01250_ ), .A2(\mreg/_04014_ ), .A3(\mreg/_01391_ ), .ZN(\mreg/_01893_ ) );
NOR4_X1 \mreg/_07781_ ( .A1(\mreg/_01890_ ), .A2(\mreg/_01891_ ), .A3(\mreg/_01892_ ), .A4(\mreg/_01893_ ), .ZN(\mreg/_01894_ ) );
NAND4_X1 \mreg/_07782_ ( .A1(\mreg/_01878_ ), .A2(\mreg/_01884_ ), .A3(\mreg/_01889_ ), .A4(\mreg/_01894_ ), .ZN(\mreg/_03918_ ) );
AND3_X1 \mreg/_07783_ ( .A1(\mreg/_01107_ ), .A2(\mreg/_01103_ ), .A3(\mreg/_04271_ ), .ZN(\mreg/_01895_ ) );
AOI221_X4 \mreg/_07784_ ( .A(\mreg/_01895_ ), .B1(\mreg/_01106_ ), .B2(\mreg/_04719_ ), .C1(\mreg/_04623_ ), .C2(\mreg/_01221_ ), .ZN(\mreg/_01896_ ) );
AND3_X1 \mreg/_07785_ ( .A1(\mreg/_01125_ ), .A2(\mreg/_04879_ ), .A3(\mreg/_01127_ ), .ZN(\mreg/_01897_ ) );
NAND3_X1 \mreg/_07786_ ( .A1(\mreg/_01117_ ), .A2(\mreg/_01103_ ), .A3(\mreg/_03951_ ), .ZN(\mreg/_01898_ ) );
INV_X1 \mreg/_07787_ ( .A(\mreg/_03983_ ), .ZN(\mreg/_01899_ ) );
OAI21_X1 \mreg/_07788_ ( .A(\mreg/_01898_ ), .B1(\mreg/_01899_ ), .B2(\mreg/_01396_ ), .ZN(\mreg/_01900_ ) );
AOI211_X4 \mreg/_07789_ ( .A(\mreg/_01897_ ), .B(\mreg/_01900_ ), .C1(\mreg/_04911_ ), .C2(\mreg/_01363_ ), .ZN(\mreg/_01901_ ) );
AND3_X1 \mreg/_07790_ ( .A1(\mreg/_01092_ ), .A2(\mreg/_01114_ ), .A3(\mreg/_04815_ ), .ZN(\mreg/_01902_ ) );
AND3_X1 \mreg/_07791_ ( .A1(\mreg/_01380_ ), .A2(\mreg/_01118_ ), .A3(\mreg/_04847_ ), .ZN(\mreg/_01903_ ) );
AND3_X1 \mreg/_07792_ ( .A1(\mreg/_01058_ ), .A2(\mreg/_01122_ ), .A3(\mreg/_04783_ ), .ZN(\mreg/_01904_ ) );
AND3_X1 \mreg/_07793_ ( .A1(\mreg/_01126_ ), .A2(\mreg/_04751_ ), .A3(\mreg/_01086_ ), .ZN(\mreg/_01905_ ) );
NOR4_X1 \mreg/_07794_ ( .A1(\mreg/_01902_ ), .A2(\mreg/_01903_ ), .A3(\mreg/_01904_ ), .A4(\mreg/_01905_ ), .ZN(\mreg/_01906_ ) );
NAND3_X1 \mreg/_07795_ ( .A1(\mreg/_01291_ ), .A2(\mreg/_04015_ ), .A3(\mreg/_01151_ ), .ZN(\mreg/_01907_ ) );
NAND3_X1 \mreg/_07796_ ( .A1(\mreg/_01143_ ), .A2(\mreg/_01114_ ), .A3(\mreg/_04079_ ), .ZN(\mreg/_01908_ ) );
NAND3_X1 \mreg/_07797_ ( .A1(\mreg/_01148_ ), .A2(\mreg/_01114_ ), .A3(\mreg/_04047_ ), .ZN(\mreg/_01909_ ) );
NAND3_X1 \mreg/_07798_ ( .A1(\mreg/_01140_ ), .A2(\mreg/_01144_ ), .A3(\mreg/_04111_ ), .ZN(\mreg/_01910_ ) );
AND4_X1 \mreg/_07799_ ( .A1(\mreg/_01907_ ), .A2(\mreg/_01908_ ), .A3(\mreg/_01909_ ), .A4(\mreg/_01910_ ), .ZN(\mreg/_01911_ ) );
AND4_X1 \mreg/_07800_ ( .A1(\mreg/_01896_ ), .A2(\mreg/_01901_ ), .A3(\mreg/_01906_ ), .A4(\mreg/_01911_ ), .ZN(\mreg/_01912_ ) );
NAND3_X1 \mreg/_07801_ ( .A1(\mreg/_01084_ ), .A2(\mreg/_04559_ ), .A3(\mreg/_01299_ ), .ZN(\mreg/_01913_ ) );
NAND4_X1 \mreg/_07802_ ( .A1(\mreg/_01365_ ), .A2(\mreg/_01366_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04495_ ), .ZN(\mreg/_01914_ ) );
INV_X1 \mreg/_07803_ ( .A(\mreg/_04527_ ), .ZN(\mreg/_01915_ ) );
OAI21_X1 \mreg/_07804_ ( .A(\mreg/_01914_ ), .B1(\mreg/_01190_ ), .B2(\mreg/_01915_ ), .ZN(\mreg/_01916_ ) );
AOI221_X4 \mreg/_07805_ ( .A(\mreg/_01916_ ), .B1(\mreg/_04463_ ), .B2(\mreg/_01195_ ), .C1(\mreg/_04431_ ), .C2(\mreg/_01660_ ), .ZN(\mreg/_01917_ ) );
NAND3_X1 \mreg/_07806_ ( .A1(\mreg/_01305_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04591_ ), .ZN(\mreg/_01918_ ) );
AND3_X1 \mreg/_07807_ ( .A1(\mreg/_01142_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04655_ ), .ZN(\mreg/_01919_ ) );
INV_X1 \mreg/_07808_ ( .A(\mreg/_00048_ ), .ZN(\mreg/_01920_ ) );
AOI21_X1 \mreg/_07809_ ( .A(\mreg/_01919_ ), .B1(\mreg/_01920_ ), .B2(\mreg/_01173_ ), .ZN(\mreg/_01921_ ) );
AND4_X1 \mreg/_07810_ ( .A1(\mreg/_01913_ ), .A2(\mreg/_01917_ ), .A3(\mreg/_01918_ ), .A4(\mreg/_01921_ ), .ZN(\mreg/_01922_ ) );
NAND4_X1 \mreg/_07811_ ( .A1(\mreg/_01667_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04207_ ), .A4(\mreg/_01212_ ), .ZN(\mreg/_01923_ ) );
INV_X1 \mreg/_07812_ ( .A(\mreg/_04239_ ), .ZN(\mreg/_01924_ ) );
OAI21_X1 \mreg/_07813_ ( .A(\mreg/_01923_ ), .B1(\mreg/_01069_ ), .B2(\mreg/_01924_ ), .ZN(\mreg/_01925_ ) );
AOI221_X4 \mreg/_07814_ ( .A(\mreg/_01925_ ), .B1(\mreg/_04175_ ), .B2(\mreg/_01075_ ), .C1(\mreg/_04143_ ), .C2(\mreg/_01080_ ), .ZN(\mreg/_01926_ ) );
NAND3_X1 \mreg/_07815_ ( .A1(\mreg/_01091_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04367_ ), .ZN(\mreg/_01927_ ) );
NAND3_X1 \mreg/_07816_ ( .A1(\mreg/_01380_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04399_ ), .ZN(\mreg/_01928_ ) );
NAND2_X1 \mreg/_07817_ ( .A1(\mreg/_01927_ ), .A2(\mreg/_01928_ ), .ZN(\mreg/_01929_ ) );
AOI221_X4 \mreg/_07818_ ( .A(\mreg/_01929_ ), .B1(\mreg/_04335_ ), .B2(\mreg/_01205_ ), .C1(\mreg/_04303_ ), .C2(\mreg/_01207_ ), .ZN(\mreg/_01930_ ) );
NAND4_X1 \mreg/_07819_ ( .A1(\mreg/_01912_ ), .A2(\mreg/_01922_ ), .A3(\mreg/_01926_ ), .A4(\mreg/_01930_ ), .ZN(\mreg/_03919_ ) );
NAND3_X1 \mreg/_07820_ ( .A1(\mreg/_01147_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04592_ ), .ZN(\mreg/_01931_ ) );
NAND3_X1 \mreg/_07821_ ( .A1(\mreg/_01255_ ), .A2(\mreg/_04560_ ), .A3(\mreg/_01150_ ), .ZN(\mreg/_01932_ ) );
NAND2_X1 \mreg/_07822_ ( .A1(\mreg/_01931_ ), .A2(\mreg/_01932_ ), .ZN(\mreg/_01933_ ) );
INV_X1 \mreg/_07823_ ( .A(\mreg/_00049_ ), .ZN(\mreg/_01934_ ) );
AOI221_X1 \mreg/_07824_ ( .A(\mreg/_01933_ ), .B1(\mreg/_01934_ ), .B2(\mreg/_01173_ ), .C1(\mreg/_04656_ ), .C2(\mreg/_01175_ ), .ZN(\mreg/_01935_ ) );
NAND4_X1 \mreg/_07825_ ( .A1(\mreg/_01318_ ), .A2(\mreg/_01453_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04496_ ), .ZN(\mreg/_01936_ ) );
INV_X1 \mreg/_07826_ ( .A(\mreg/_04528_ ), .ZN(\mreg/_01937_ ) );
OAI21_X1 \mreg/_07827_ ( .A(\mreg/_01936_ ), .B1(\mreg/_01678_ ), .B2(\mreg/_01937_ ), .ZN(\mreg/_01938_ ) );
AOI221_X4 \mreg/_07828_ ( .A(\mreg/_01938_ ), .B1(\mreg/_04464_ ), .B2(\mreg/_01412_ ), .C1(\mreg/_04432_ ), .C2(\mreg/_01198_ ), .ZN(\mreg/_01939_ ) );
NAND3_X1 \mreg/_07829_ ( .A1(\mreg/_01323_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04368_ ), .ZN(\mreg/_01940_ ) );
NAND3_X1 \mreg/_07830_ ( .A1(\mreg/_01496_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04400_ ), .ZN(\mreg/_01941_ ) );
NAND2_X1 \mreg/_07831_ ( .A1(\mreg/_01940_ ), .A2(\mreg/_01941_ ), .ZN(\mreg/_01942_ ) );
AOI221_X4 \mreg/_07832_ ( .A(\mreg/_01942_ ), .B1(\mreg/_04336_ ), .B2(\mreg/_01611_ ), .C1(\mreg/_04304_ ), .C2(\mreg/_01499_ ), .ZN(\mreg/_01943_ ) );
NAND4_X1 \mreg/_07833_ ( .A1(\mreg/_01501_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04208_ ), .A4(\mreg/_01372_ ), .ZN(\mreg/_01944_ ) );
INV_X1 \mreg/_07834_ ( .A(\mreg/_04240_ ), .ZN(\mreg/_01945_ ) );
OAI21_X1 \mreg/_07835_ ( .A(\mreg/_01944_ ), .B1(\mreg/_01374_ ), .B2(\mreg/_01945_ ), .ZN(\mreg/_01946_ ) );
AOI221_X4 \mreg/_07836_ ( .A(\mreg/_01946_ ), .B1(\mreg/_04176_ ), .B2(\mreg/_01465_ ), .C1(\mreg/_04144_ ), .C2(\mreg/_01505_ ), .ZN(\mreg/_01947_ ) );
AND4_X4 \mreg/_07837_ ( .A1(\mreg/_01935_ ), .A2(\mreg/_01939_ ), .A3(\mreg/_01943_ ), .A4(\mreg/_01947_ ), .ZN(\mreg/_01948_ ) );
NAND3_X1 \mreg/_07838_ ( .A1(\mreg/_01275_ ), .A2(\mreg/_01277_ ), .A3(\mreg/_04816_ ), .ZN(\mreg/_01949_ ) );
AOI22_X1 \mreg/_07839_ ( .A1(\mreg/_01284_ ), .A2(\mreg/_04784_ ), .B1(\mreg/_04752_ ), .B2(\mreg/_01230_ ), .ZN(\mreg/_01950_ ) );
NAND3_X1 \mreg/_07840_ ( .A1(\mreg/_01281_ ), .A2(\mreg/_01302_ ), .A3(\mreg/_04848_ ), .ZN(\mreg/_01951_ ) );
NAND3_X1 \mreg/_07841_ ( .A1(\mreg/_01621_ ), .A2(\mreg/_01622_ ), .A3(\mreg/_04272_ ), .ZN(\mreg/_01952_ ) );
NAND3_X1 \mreg/_07842_ ( .A1(\mreg/_01386_ ), .A2(\mreg/_01622_ ), .A3(\mreg/_04624_ ), .ZN(\mreg/_01953_ ) );
NAND3_X1 \mreg/_07843_ ( .A1(\mreg/_01067_ ), .A2(\mreg/_01130_ ), .A3(\mreg/_04720_ ), .ZN(\mreg/_01954_ ) );
AND3_X1 \mreg/_07844_ ( .A1(\mreg/_01952_ ), .A2(\mreg/_01953_ ), .A3(\mreg/_01954_ ), .ZN(\mreg/_01955_ ) );
AND4_X1 \mreg/_07845_ ( .A1(\mreg/_01949_ ), .A2(\mreg/_01950_ ), .A3(\mreg/_01951_ ), .A4(\mreg/_01955_ ), .ZN(\mreg/_01956_ ) );
AND3_X1 \mreg/_07846_ ( .A1(\mreg/_01112_ ), .A2(\mreg/_01217_ ), .A3(\mreg/_03984_ ), .ZN(\mreg/_01957_ ) );
NAND3_X1 \mreg/_07847_ ( .A1(\mreg/_01121_ ), .A2(\mreg/_01144_ ), .A3(\mreg/_04912_ ), .ZN(\mreg/_01958_ ) );
NAND3_X1 \mreg/_07848_ ( .A1(\mreg/_01338_ ), .A2(\mreg/_01162_ ), .A3(\mreg/_04880_ ), .ZN(\mreg/_01959_ ) );
NAND2_X1 \mreg/_07849_ ( .A1(\mreg/_01958_ ), .A2(\mreg/_01959_ ), .ZN(\mreg/_01960_ ) );
AOI211_X4 \mreg/_07850_ ( .A(\mreg/_01957_ ), .B(\mreg/_01960_ ), .C1(\mreg/_03952_ ), .C2(\mreg/_01361_ ), .ZN(\mreg/_01961_ ) );
AND3_X1 \mreg/_07851_ ( .A1(\mreg/_01232_ ), .A2(\mreg/_01233_ ), .A3(\mreg/_04080_ ), .ZN(\mreg/_01962_ ) );
AND3_X1 \mreg/_07852_ ( .A1(\mreg/_01304_ ), .A2(\mreg/_01384_ ), .A3(\mreg/_04048_ ), .ZN(\mreg/_01963_ ) );
AND3_X1 \mreg/_07853_ ( .A1(\mreg/_01238_ ), .A2(\mreg/_01248_ ), .A3(\mreg/_04112_ ), .ZN(\mreg/_01964_ ) );
AND3_X1 \mreg/_07854_ ( .A1(\mreg/_01250_ ), .A2(\mreg/_04016_ ), .A3(\mreg/_01391_ ), .ZN(\mreg/_01965_ ) );
NOR4_X1 \mreg/_07855_ ( .A1(\mreg/_01962_ ), .A2(\mreg/_01963_ ), .A3(\mreg/_01964_ ), .A4(\mreg/_01965_ ), .ZN(\mreg/_01966_ ) );
NAND4_X1 \mreg/_07856_ ( .A1(\mreg/_01948_ ), .A2(\mreg/_01956_ ), .A3(\mreg/_01961_ ), .A4(\mreg/_01966_ ), .ZN(\mreg/_03920_ ) );
NAND3_X1 \mreg/_07857_ ( .A1(\mreg/_01083_ ), .A2(\mreg/_04562_ ), .A3(\mreg/_01597_ ), .ZN(\mreg/_01967_ ) );
NAND3_X1 \mreg/_07858_ ( .A1(\mreg/_01180_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04658_ ), .ZN(\mreg/_01968_ ) );
NAND3_X1 \mreg/_07859_ ( .A1(\mreg/_01182_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04594_ ), .ZN(\mreg/_01969_ ) );
INV_X1 \mreg/_07860_ ( .A(\mreg/_00050_ ), .ZN(\mreg/_01970_ ) );
NAND3_X1 \mreg/_07861_ ( .A1(\mreg/_01184_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_01970_ ), .ZN(\mreg/_01971_ ) );
AND4_X1 \mreg/_07862_ ( .A1(\mreg/_01967_ ), .A2(\mreg/_01968_ ), .A3(\mreg/_01969_ ), .A4(\mreg/_01971_ ), .ZN(\mreg/_01972_ ) );
NAND4_X1 \mreg/_07863_ ( .A1(\mreg/_01269_ ), .A2(\mreg/_01453_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04498_ ), .ZN(\mreg/_01973_ ) );
INV_X1 \mreg/_07864_ ( .A(\mreg/_04530_ ), .ZN(\mreg/_01974_ ) );
OAI21_X1 \mreg/_07865_ ( .A(\mreg/_01973_ ), .B1(\mreg/_01678_ ), .B2(\mreg/_01974_ ), .ZN(\mreg/_01975_ ) );
AOI221_X4 \mreg/_07866_ ( .A(\mreg/_01975_ ), .B1(\mreg/_04466_ ), .B2(\mreg/_01412_ ), .C1(\mreg/_04434_ ), .C2(\mreg/_01660_ ), .ZN(\mreg/_01976_ ) );
NAND3_X1 \mreg/_07867_ ( .A1(\mreg/_01323_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04370_ ), .ZN(\mreg/_01977_ ) );
NAND3_X1 \mreg/_07868_ ( .A1(\mreg/_01496_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04402_ ), .ZN(\mreg/_01978_ ) );
NAND2_X1 \mreg/_07869_ ( .A1(\mreg/_01977_ ), .A2(\mreg/_01978_ ), .ZN(\mreg/_01979_ ) );
AOI221_X4 \mreg/_07870_ ( .A(\mreg/_01979_ ), .B1(\mreg/_04338_ ), .B2(\mreg/_01611_ ), .C1(\mreg/_04306_ ), .C2(\mreg/_01499_ ), .ZN(\mreg/_01980_ ) );
BUF_X4 \mreg/_07871_ ( .A(\mreg/_01212_ ), .Z(\mreg/_01981_ ) );
NAND3_X1 \mreg/_07872_ ( .A1(\mreg/_01082_ ), .A2(\mreg/_04146_ ), .A3(\mreg/_01981_ ), .ZN(\mreg/_01982_ ) );
NAND3_X1 \mreg/_07873_ ( .A1(\mreg/_01621_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04178_ ), .ZN(\mreg/_01983_ ) );
NAND4_X1 \mreg/_07874_ ( .A1(\mreg/_01667_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04210_ ), .A4(\mreg/_01981_ ), .ZN(\mreg/_01984_ ) );
NAND4_X1 \mreg/_07875_ ( .A1(\mreg/_01211_ ), .A2(\mreg/_01981_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04242_ ), .ZN(\mreg/_01985_ ) );
AND4_X1 \mreg/_07876_ ( .A1(\mreg/_01982_ ), .A2(\mreg/_01983_ ), .A3(\mreg/_01984_ ), .A4(\mreg/_01985_ ), .ZN(\mreg/_01986_ ) );
AND4_X4 \mreg/_07877_ ( .A1(\mreg/_01972_ ), .A2(\mreg/_01976_ ), .A3(\mreg/_01980_ ), .A4(\mreg/_01986_ ), .ZN(\mreg/_01987_ ) );
NAND3_X1 \mreg/_07878_ ( .A1(\mreg/_01059_ ), .A2(\mreg/_01277_ ), .A3(\mreg/_04786_ ), .ZN(\mreg/_01988_ ) );
AND3_X1 \mreg/_07879_ ( .A1(\mreg/_01064_ ), .A2(\mreg/_01357_ ), .A3(\mreg/_04626_ ), .ZN(\mreg/_01989_ ) );
AOI221_X4 \mreg/_07880_ ( .A(\mreg/_01989_ ), .B1(\mreg/_01106_ ), .B2(\mreg/_04722_ ), .C1(\mreg/_04274_ ), .C2(\mreg/_01110_ ), .ZN(\mreg/_01990_ ) );
NAND3_X1 \mreg/_07881_ ( .A1(\mreg/_01298_ ), .A2(\mreg/_01087_ ), .A3(\mreg/_04754_ ), .ZN(\mreg/_01991_ ) );
AND3_X1 \mreg/_07882_ ( .A1(\mreg/_01098_ ), .A2(\mreg/_01133_ ), .A3(\mreg/_04850_ ), .ZN(\mreg/_01992_ ) );
AOI21_X1 \mreg/_07883_ ( .A(\mreg/_01992_ ), .B1(\mreg/_04818_ ), .B2(\mreg/_01431_ ), .ZN(\mreg/_01993_ ) );
AND4_X1 \mreg/_07884_ ( .A1(\mreg/_01988_ ), .A2(\mreg/_01990_ ), .A3(\mreg/_01991_ ), .A4(\mreg/_01993_ ), .ZN(\mreg/_01994_ ) );
NAND3_X1 \mreg/_07885_ ( .A1(\mreg/_01156_ ), .A2(\mreg/_01436_ ), .A3(\mreg/_04914_ ), .ZN(\mreg/_01995_ ) );
NAND3_X1 \mreg/_07886_ ( .A1(\mreg/_01159_ ), .A2(\mreg/_01289_ ), .A3(\mreg/_03954_ ), .ZN(\mreg/_01996_ ) );
NAND3_X1 \mreg/_07887_ ( .A1(\mreg/_01292_ ), .A2(\mreg/_01293_ ), .A3(\mreg/_04882_ ), .ZN(\mreg/_01997_ ) );
NAND3_X1 \mreg/_07888_ ( .A1(\mreg/_01165_ ), .A2(\mreg/_01477_ ), .A3(\mreg/_03986_ ), .ZN(\mreg/_01998_ ) );
AND4_X1 \mreg/_07889_ ( .A1(\mreg/_01995_ ), .A2(\mreg/_01996_ ), .A3(\mreg/_01997_ ), .A4(\mreg/_01998_ ), .ZN(\mreg/_01999_ ) );
NAND3_X1 \mreg/_07890_ ( .A1(\mreg/_01298_ ), .A2(\mreg/_04018_ ), .A3(\mreg/_01299_ ), .ZN(\mreg/_02000_ ) );
NAND3_X1 \mreg/_07891_ ( .A1(\mreg/_01301_ ), .A2(\mreg/_01302_ ), .A3(\mreg/_04082_ ), .ZN(\mreg/_02001_ ) );
NAND3_X1 \mreg/_07892_ ( .A1(\mreg/_01305_ ), .A2(\mreg/_01295_ ), .A3(\mreg/_04050_ ), .ZN(\mreg/_02002_ ) );
NAND3_X1 \mreg/_07893_ ( .A1(\mreg/_01308_ ), .A2(\mreg/_01309_ ), .A3(\mreg/_04114_ ), .ZN(\mreg/_02003_ ) );
AND4_X1 \mreg/_07894_ ( .A1(\mreg/_02000_ ), .A2(\mreg/_02001_ ), .A3(\mreg/_02002_ ), .A4(\mreg/_02003_ ), .ZN(\mreg/_02004_ ) );
NAND4_X1 \mreg/_07895_ ( .A1(\mreg/_01987_ ), .A2(\mreg/_01994_ ), .A3(\mreg/_01999_ ), .A4(\mreg/_02004_ ), .ZN(\mreg/_03922_ ) );
NAND3_X1 \mreg/_07896_ ( .A1(\mreg/_01083_ ), .A2(\mreg/_04563_ ), .A3(\mreg/_01597_ ), .ZN(\mreg/_02005_ ) );
NAND3_X1 \mreg/_07897_ ( .A1(\mreg/_01180_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04659_ ), .ZN(\mreg/_02006_ ) );
NAND3_X1 \mreg/_07898_ ( .A1(\mreg/_01182_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04595_ ), .ZN(\mreg/_02007_ ) );
INV_X1 \mreg/_07899_ ( .A(\mreg/_00051_ ), .ZN(\mreg/_02008_ ) );
NAND3_X1 \mreg/_07900_ ( .A1(\mreg/_01184_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_02008_ ), .ZN(\mreg/_02009_ ) );
AND4_X1 \mreg/_07901_ ( .A1(\mreg/_02005_ ), .A2(\mreg/_02006_ ), .A3(\mreg/_02007_ ), .A4(\mreg/_02009_ ), .ZN(\mreg/_02010_ ) );
NAND4_X1 \mreg/_07902_ ( .A1(\mreg/_01269_ ), .A2(\mreg/_01453_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04499_ ), .ZN(\mreg/_02011_ ) );
INV_X1 \mreg/_07903_ ( .A(\mreg/_04531_ ), .ZN(\mreg/_02012_ ) );
OAI21_X1 \mreg/_07904_ ( .A(\mreg/_02011_ ), .B1(\mreg/_01678_ ), .B2(\mreg/_02012_ ), .ZN(\mreg/_02013_ ) );
AOI221_X4 \mreg/_07905_ ( .A(\mreg/_02013_ ), .B1(\mreg/_04467_ ), .B2(\mreg/_01412_ ), .C1(\mreg/_04435_ ), .C2(\mreg/_01660_ ), .ZN(\mreg/_02014_ ) );
NAND3_X1 \mreg/_07906_ ( .A1(\mreg/_01323_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04371_ ), .ZN(\mreg/_02015_ ) );
NAND3_X1 \mreg/_07907_ ( .A1(\mreg/_01496_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04403_ ), .ZN(\mreg/_02016_ ) );
NAND2_X1 \mreg/_07908_ ( .A1(\mreg/_02015_ ), .A2(\mreg/_02016_ ), .ZN(\mreg/_02017_ ) );
AOI221_X4 \mreg/_07909_ ( .A(\mreg/_02017_ ), .B1(\mreg/_04339_ ), .B2(\mreg/_01611_ ), .C1(\mreg/_04307_ ), .C2(\mreg/_01499_ ), .ZN(\mreg/_02018_ ) );
NAND4_X1 \mreg/_07910_ ( .A1(\mreg/_01188_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04211_ ), .A4(\mreg/_01209_ ), .ZN(\mreg/_02019_ ) );
NAND4_X1 \mreg/_07911_ ( .A1(\mreg/_01211_ ), .A2(\mreg/_01209_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04243_ ), .ZN(\mreg/_02020_ ) );
NAND2_X1 \mreg/_07912_ ( .A1(\mreg/_02019_ ), .A2(\mreg/_02020_ ), .ZN(\mreg/_02021_ ) );
AOI221_X4 \mreg/_07913_ ( .A(\mreg/_02021_ ), .B1(\mreg/_04179_ ), .B2(\mreg/_01465_ ), .C1(\mreg/_04147_ ), .C2(\mreg/_01505_ ), .ZN(\mreg/_02022_ ) );
AND4_X2 \mreg/_07914_ ( .A1(\mreg/_02010_ ), .A2(\mreg/_02014_ ), .A3(\mreg/_02018_ ), .A4(\mreg/_02022_ ), .ZN(\mreg/_02023_ ) );
NAND3_X1 \mreg/_07915_ ( .A1(\mreg/_01383_ ), .A2(\mreg/_01277_ ), .A3(\mreg/_04275_ ), .ZN(\mreg/_02024_ ) );
AND3_X1 \mreg/_07916_ ( .A1(\mreg/_01098_ ), .A2(\mreg/_01144_ ), .A3(\mreg/_04851_ ), .ZN(\mreg/_02025_ ) );
AOI21_X1 \mreg/_07917_ ( .A(\mreg/_02025_ ), .B1(\mreg/_04819_ ), .B2(\mreg/_01431_ ), .ZN(\mreg/_02026_ ) );
AOI22_X1 \mreg/_07918_ ( .A1(\mreg/_04627_ ), .A2(\mreg/_01222_ ), .B1(\mreg/_01219_ ), .B2(\mreg/_04723_ ), .ZN(\mreg/_02027_ ) );
AOI22_X1 \mreg/_07919_ ( .A1(\mreg/_01284_ ), .A2(\mreg/_04787_ ), .B1(\mreg/_04755_ ), .B2(\mreg/_01230_ ), .ZN(\mreg/_02028_ ) );
AND4_X1 \mreg/_07920_ ( .A1(\mreg/_02024_ ), .A2(\mreg/_02026_ ), .A3(\mreg/_02027_ ), .A4(\mreg/_02028_ ), .ZN(\mreg/_02029_ ) );
NAND3_X1 \mreg/_07921_ ( .A1(\mreg/_01156_ ), .A2(\mreg/_01436_ ), .A3(\mreg/_04915_ ), .ZN(\mreg/_02030_ ) );
NAND3_X1 \mreg/_07922_ ( .A1(\mreg/_01159_ ), .A2(\mreg/_01289_ ), .A3(\mreg/_03955_ ), .ZN(\mreg/_02031_ ) );
NAND3_X1 \mreg/_07923_ ( .A1(\mreg/_01292_ ), .A2(\mreg/_01293_ ), .A3(\mreg/_04883_ ), .ZN(\mreg/_02032_ ) );
NAND3_X1 \mreg/_07924_ ( .A1(\mreg/_01165_ ), .A2(\mreg/_01477_ ), .A3(\mreg/_03987_ ), .ZN(\mreg/_02033_ ) );
AND4_X1 \mreg/_07925_ ( .A1(\mreg/_02030_ ), .A2(\mreg/_02031_ ), .A3(\mreg/_02032_ ), .A4(\mreg/_02033_ ), .ZN(\mreg/_02034_ ) );
NAND3_X1 \mreg/_07926_ ( .A1(\mreg/_01298_ ), .A2(\mreg/_04019_ ), .A3(\mreg/_01299_ ), .ZN(\mreg/_02035_ ) );
NAND3_X1 \mreg/_07927_ ( .A1(\mreg/_01301_ ), .A2(\mreg/_01302_ ), .A3(\mreg/_04083_ ), .ZN(\mreg/_02036_ ) );
NAND3_X1 \mreg/_07928_ ( .A1(\mreg/_01235_ ), .A2(\mreg/_01295_ ), .A3(\mreg/_04051_ ), .ZN(\mreg/_02037_ ) );
NAND3_X1 \mreg/_07929_ ( .A1(\mreg/_01308_ ), .A2(\mreg/_01309_ ), .A3(\mreg/_04115_ ), .ZN(\mreg/_02038_ ) );
AND4_X1 \mreg/_07930_ ( .A1(\mreg/_02035_ ), .A2(\mreg/_02036_ ), .A3(\mreg/_02037_ ), .A4(\mreg/_02038_ ), .ZN(\mreg/_02039_ ) );
NAND4_X1 \mreg/_07931_ ( .A1(\mreg/_02023_ ), .A2(\mreg/_02029_ ), .A3(\mreg/_02034_ ), .A4(\mreg/_02039_ ), .ZN(\mreg/_03923_ ) );
NAND3_X1 \mreg/_07932_ ( .A1(\mreg/_01083_ ), .A2(\mreg/_04564_ ), .A3(\mreg/_01597_ ), .ZN(\mreg/_02040_ ) );
NAND3_X1 \mreg/_07933_ ( .A1(\mreg/_01143_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04660_ ), .ZN(\mreg/_02041_ ) );
NAND3_X1 \mreg/_07934_ ( .A1(\mreg/_01182_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04596_ ), .ZN(\mreg/_02042_ ) );
INV_X1 \mreg/_07935_ ( .A(\mreg/_00052_ ), .ZN(\mreg/_02043_ ) );
NAND3_X1 \mreg/_07936_ ( .A1(\mreg/_01140_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_02043_ ), .ZN(\mreg/_02044_ ) );
AND4_X1 \mreg/_07937_ ( .A1(\mreg/_02040_ ), .A2(\mreg/_02041_ ), .A3(\mreg/_02042_ ), .A4(\mreg/_02044_ ), .ZN(\mreg/_02045_ ) );
NAND4_X1 \mreg/_07938_ ( .A1(\mreg/_01269_ ), .A2(\mreg/_01366_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04500_ ), .ZN(\mreg/_02046_ ) );
INV_X1 \mreg/_07939_ ( .A(\mreg/_04532_ ), .ZN(\mreg/_02047_ ) );
OAI21_X1 \mreg/_07940_ ( .A(\mreg/_02046_ ), .B1(\mreg/_01678_ ), .B2(\mreg/_02047_ ), .ZN(\mreg/_02048_ ) );
AOI221_X4 \mreg/_07941_ ( .A(\mreg/_02048_ ), .B1(\mreg/_04468_ ), .B2(\mreg/_01195_ ), .C1(\mreg/_04436_ ), .C2(\mreg/_01660_ ), .ZN(\mreg/_02049_ ) );
NAND3_X1 \mreg/_07942_ ( .A1(\mreg/_01398_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04372_ ), .ZN(\mreg/_02050_ ) );
NAND3_X1 \mreg/_07943_ ( .A1(\mreg/_01496_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04404_ ), .ZN(\mreg/_02051_ ) );
NAND2_X1 \mreg/_07944_ ( .A1(\mreg/_02050_ ), .A2(\mreg/_02051_ ), .ZN(\mreg/_02052_ ) );
AOI221_X4 \mreg/_07945_ ( .A(\mreg/_02052_ ), .B1(\mreg/_04340_ ), .B2(\mreg/_01611_ ), .C1(\mreg/_04308_ ), .C2(\mreg/_01499_ ), .ZN(\mreg/_02053_ ) );
NAND3_X1 \mreg/_07946_ ( .A1(\mreg/_01082_ ), .A2(\mreg/_04148_ ), .A3(\mreg/_01981_ ), .ZN(\mreg/_02054_ ) );
NAND3_X1 \mreg/_07947_ ( .A1(\mreg/_01621_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04180_ ), .ZN(\mreg/_02055_ ) );
NAND4_X1 \mreg/_07948_ ( .A1(\mreg/_01667_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04212_ ), .A4(\mreg/_01212_ ), .ZN(\mreg/_02056_ ) );
NAND4_X1 \mreg/_07949_ ( .A1(\mreg/_01211_ ), .A2(\mreg/_01981_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04244_ ), .ZN(\mreg/_02057_ ) );
AND4_X1 \mreg/_07950_ ( .A1(\mreg/_02054_ ), .A2(\mreg/_02055_ ), .A3(\mreg/_02056_ ), .A4(\mreg/_02057_ ), .ZN(\mreg/_02058_ ) );
AND4_X2 \mreg/_07951_ ( .A1(\mreg/_02045_ ), .A2(\mreg/_02049_ ), .A3(\mreg/_02053_ ), .A4(\mreg/_02058_ ), .ZN(\mreg/_02059_ ) );
AND3_X1 \mreg/_07952_ ( .A1(\mreg/_01107_ ), .A2(\mreg/_01217_ ), .A3(\mreg/_04276_ ), .ZN(\mreg/_02060_ ) );
AOI221_X4 \mreg/_07953_ ( .A(\mreg/_02060_ ), .B1(\mreg/_01219_ ), .B2(\mreg/_04724_ ), .C1(\mreg/_04628_ ), .C2(\mreg/_01222_ ), .ZN(\mreg/_02061_ ) );
NAND3_X1 \mreg/_07954_ ( .A1(\mreg/_01059_ ), .A2(\mreg/_01436_ ), .A3(\mreg/_04788_ ), .ZN(\mreg/_02062_ ) );
NAND3_X1 \mreg/_07955_ ( .A1(\mreg/_01092_ ), .A2(\mreg/_01282_ ), .A3(\mreg/_04820_ ), .ZN(\mreg/_02063_ ) );
NAND3_X1 \mreg/_07956_ ( .A1(\mreg/_01381_ ), .A2(\mreg/_01306_ ), .A3(\mreg/_04852_ ), .ZN(\mreg/_02064_ ) );
NAND3_X1 \mreg/_07957_ ( .A1(\mreg/_01339_ ), .A2(\mreg/_01087_ ), .A3(\mreg/_04756_ ), .ZN(\mreg/_02065_ ) );
AND4_X1 \mreg/_07958_ ( .A1(\mreg/_02062_ ), .A2(\mreg/_02063_ ), .A3(\mreg/_02064_ ), .A4(\mreg/_02065_ ), .ZN(\mreg/_02066_ ) );
NAND3_X1 \mreg/_07959_ ( .A1(\mreg/_01232_ ), .A2(\mreg/_01233_ ), .A3(\mreg/_04084_ ), .ZN(\mreg/_02067_ ) );
NAND3_X1 \mreg/_07960_ ( .A1(\mreg/_01235_ ), .A2(\mreg/_01236_ ), .A3(\mreg/_04052_ ), .ZN(\mreg/_02068_ ) );
NAND3_X1 \mreg/_07961_ ( .A1(\mreg/_01238_ ), .A2(\mreg/_01239_ ), .A3(\mreg/_04116_ ), .ZN(\mreg/_02069_ ) );
NAND3_X1 \mreg/_07962_ ( .A1(\mreg/_01241_ ), .A2(\mreg/_04020_ ), .A3(\mreg/_01242_ ), .ZN(\mreg/_02070_ ) );
NAND4_X1 \mreg/_07963_ ( .A1(\mreg/_02067_ ), .A2(\mreg/_02068_ ), .A3(\mreg/_02069_ ), .A4(\mreg/_02070_ ), .ZN(\mreg/_02071_ ) );
NAND3_X1 \mreg/_07964_ ( .A1(\mreg/_01158_ ), .A2(\mreg/_01236_ ), .A3(\mreg/_03956_ ), .ZN(\mreg/_02072_ ) );
NAND3_X1 \mreg/_07965_ ( .A1(\mreg/_01113_ ), .A2(\mreg/_01236_ ), .A3(\mreg/_03988_ ), .ZN(\mreg/_02073_ ) );
NAND2_X1 \mreg/_07966_ ( .A1(\mreg/_02072_ ), .A2(\mreg/_02073_ ), .ZN(\mreg/_02074_ ) );
AND3_X1 \mreg/_07967_ ( .A1(\mreg/_01155_ ), .A2(\mreg/_01248_ ), .A3(\mreg/_04916_ ), .ZN(\mreg/_02075_ ) );
AND3_X1 \mreg/_07968_ ( .A1(\mreg/_01250_ ), .A2(\mreg/_04884_ ), .A3(\mreg/_01251_ ), .ZN(\mreg/_02076_ ) );
NOR4_X1 \mreg/_07969_ ( .A1(\mreg/_02071_ ), .A2(\mreg/_02074_ ), .A3(\mreg/_02075_ ), .A4(\mreg/_02076_ ), .ZN(\mreg/_02077_ ) );
NAND4_X1 \mreg/_07970_ ( .A1(\mreg/_02059_ ), .A2(\mreg/_02061_ ), .A3(\mreg/_02066_ ), .A4(\mreg/_02077_ ), .ZN(\mreg/_03924_ ) );
NAND3_X1 \mreg/_07971_ ( .A1(\mreg/_01125_ ), .A2(\mreg/_01086_ ), .A3(\mreg/_04757_ ), .ZN(\mreg/_02078_ ) );
INV_X1 \mreg/_07972_ ( .A(\mreg/_04725_ ), .ZN(\mreg/_02079_ ) );
OAI21_X1 \mreg/_07973_ ( .A(\mreg/_02078_ ), .B1(\mreg/_01786_ ), .B2(\mreg/_02079_ ), .ZN(\mreg/_02080_ ) );
AOI221_X1 \mreg/_07974_ ( .A(\mreg/_02080_ ), .B1(\mreg/_04821_ ), .B2(\mreg/_01430_ ), .C1(\mreg/_04789_ ), .C2(\mreg/_01228_ ), .ZN(\mreg/_02081_ ) );
NAND3_X1 \mreg/_07975_ ( .A1(\mreg/_01139_ ), .A2(\mreg/_01108_ ), .A3(\mreg/_04117_ ), .ZN(\mreg/_02082_ ) );
INV_X1 \mreg/_07976_ ( .A(\mreg/_04053_ ), .ZN(\mreg/_02083_ ) );
OAI21_X1 \mreg/_07977_ ( .A(\mreg/_02082_ ), .B1(\mreg/_01791_ ), .B2(\mreg/_02083_ ), .ZN(\mreg/_02084_ ) );
AOI221_X1 \mreg/_07978_ ( .A(\mreg/_02084_ ), .B1(\mreg/_03957_ ), .B2(\mreg/_01361_ ), .C1(\mreg/_04917_ ), .C2(\mreg/_01363_ ), .ZN(\mreg/_02085_ ) );
NAND4_X1 \mreg/_07979_ ( .A1(\mreg/_01365_ ), .A2(\mreg/_01116_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04501_ ), .ZN(\mreg/_02086_ ) );
INV_X1 \mreg/_07980_ ( .A(\mreg/_04533_ ), .ZN(\mreg/_02087_ ) );
OAI21_X1 \mreg/_07981_ ( .A(\mreg/_02086_ ), .B1(\mreg/_01190_ ), .B2(\mreg/_02087_ ), .ZN(\mreg/_02088_ ) );
INV_X1 \mreg/_07982_ ( .A(\mreg/_00053_ ), .ZN(\mreg/_02089_ ) );
AOI221_X1 \mreg/_07983_ ( .A(\mreg/_02088_ ), .B1(\mreg/_02089_ ), .B2(\mreg/_01172_ ), .C1(\mreg/_04661_ ), .C2(\mreg/_01174_ ), .ZN(\mreg/_02090_ ) );
NAND4_X1 \mreg/_07984_ ( .A1(\mreg/_01089_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04213_ ), .A4(\mreg/_01062_ ), .ZN(\mreg/_02091_ ) );
INV_X1 \mreg/_07985_ ( .A(\mreg/_04245_ ), .ZN(\mreg/_02092_ ) );
OAI21_X1 \mreg/_07986_ ( .A(\mreg/_02091_ ), .B1(\mreg/_01068_ ), .B2(\mreg/_02092_ ), .ZN(\mreg/_02093_ ) );
AOI221_X4 \mreg/_07987_ ( .A(\mreg/_02093_ ), .B1(\mreg/_04341_ ), .B2(\mreg/_01204_ ), .C1(\mreg/_04309_ ), .C2(\mreg/_01377_ ), .ZN(\mreg/_02094_ ) );
NAND4_X1 \mreg/_07988_ ( .A1(\mreg/_02081_ ), .A2(\mreg/_02085_ ), .A3(\mreg/_02090_ ), .A4(\mreg/_02094_ ), .ZN(\mreg/_02095_ ) );
NAND3_X1 \mreg/_07989_ ( .A1(\mreg/_01381_ ), .A2(\mreg/_01239_ ), .A3(\mreg/_04853_ ), .ZN(\mreg/_02096_ ) );
NAND3_X1 \mreg/_07990_ ( .A1(\mreg/_01621_ ), .A2(\mreg/_01384_ ), .A3(\mreg/_04277_ ), .ZN(\mreg/_02097_ ) );
NAND3_X1 \mreg/_07991_ ( .A1(\mreg/_01386_ ), .A2(\mreg/_01387_ ), .A3(\mreg/_04629_ ), .ZN(\mreg/_02098_ ) );
NAND3_X1 \mreg/_07992_ ( .A1(\mreg/_01241_ ), .A2(\mreg/_01163_ ), .A3(\mreg/_04885_ ), .ZN(\mreg/_02099_ ) );
NAND4_X1 \mreg/_07993_ ( .A1(\mreg/_02096_ ), .A2(\mreg/_02097_ ), .A3(\mreg/_02098_ ), .A4(\mreg/_02099_ ), .ZN(\mreg/_02100_ ) );
NAND3_X1 \mreg/_07994_ ( .A1(\mreg/_01291_ ), .A2(\mreg/_04021_ ), .A3(\mreg/_01391_ ), .ZN(\mreg/_02101_ ) );
INV_X1 \mreg/_07995_ ( .A(\mreg/_04085_ ), .ZN(\mreg/_02102_ ) );
INV_X1 \mreg/_07996_ ( .A(\mreg/_03989_ ), .ZN(\mreg/_02103_ ) );
OAI221_X1 \mreg/_07997_ ( .A(\mreg/_02101_ ), .B1(\mreg/_01393_ ), .B2(\mreg/_02102_ ), .C1(\mreg/_02103_ ), .C2(\mreg/_01396_ ), .ZN(\mreg/_02104_ ) );
NAND3_X1 \mreg/_07998_ ( .A1(\mreg/_01398_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04373_ ), .ZN(\mreg/_02105_ ) );
NAND3_X2 \mreg/_07999_ ( .A1(\mreg/_01096_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04405_ ), .ZN(\mreg/_02106_ ) );
NAND2_X1 \mreg/_08000_ ( .A1(\mreg/_02105_ ), .A2(\mreg/_02106_ ), .ZN(\mreg/_02107_ ) );
AOI221_X1 \mreg/_08001_ ( .A(\mreg/_02107_ ), .B1(\mreg/_04181_ ), .B2(\mreg/_01074_ ), .C1(\mreg/_04149_ ), .C2(\mreg/_01079_ ), .ZN(\mreg/_02108_ ) );
NAND3_X1 \mreg/_08002_ ( .A1(\mreg/_01177_ ), .A2(\mreg/_04565_ ), .A3(\mreg/_01391_ ), .ZN(\mreg/_02109_ ) );
NAND3_X1 \mreg/_08003_ ( .A1(\mreg/_01304_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04597_ ), .ZN(\mreg/_02110_ ) );
NAND3_X1 \mreg/_08004_ ( .A1(\mreg/_01121_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04469_ ), .ZN(\mreg/_02111_ ) );
NAND3_X1 \mreg/_08005_ ( .A1(\mreg/_01082_ ), .A2(\mreg/_04437_ ), .A3(\mreg/_01162_ ), .ZN(\mreg/_02112_ ) );
AND2_X1 \mreg/_08006_ ( .A1(\mreg/_02111_ ), .A2(\mreg/_02112_ ), .ZN(\mreg/_02113_ ) );
NAND4_X1 \mreg/_08007_ ( .A1(\mreg/_02108_ ), .A2(\mreg/_02109_ ), .A3(\mreg/_02110_ ), .A4(\mreg/_02113_ ), .ZN(\mreg/_02114_ ) );
OR4_X2 \mreg/_08008_ ( .A1(\mreg/_02095_ ), .A2(\mreg/_02100_ ), .A3(\mreg/_02104_ ), .A4(\mreg/_02114_ ), .ZN(\mreg/_03925_ ) );
NAND3_X1 \mreg/_08009_ ( .A1(\mreg/_01147_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04598_ ), .ZN(\mreg/_02115_ ) );
NAND3_X1 \mreg/_08010_ ( .A1(\mreg/_01255_ ), .A2(\mreg/_04566_ ), .A3(\mreg/_01150_ ), .ZN(\mreg/_02116_ ) );
NAND2_X1 \mreg/_08011_ ( .A1(\mreg/_02115_ ), .A2(\mreg/_02116_ ), .ZN(\mreg/_02117_ ) );
INV_X1 \mreg/_08012_ ( .A(\mreg/_00054_ ), .ZN(\mreg/_02118_ ) );
AOI221_X1 \mreg/_08013_ ( .A(\mreg/_02117_ ), .B1(\mreg/_02118_ ), .B2(\mreg/_01173_ ), .C1(\mreg/_04662_ ), .C2(\mreg/_01175_ ), .ZN(\mreg/_02119_ ) );
NAND4_X1 \mreg/_08014_ ( .A1(\mreg/_01269_ ), .A2(\mreg/_01366_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04502_ ), .ZN(\mreg/_02120_ ) );
INV_X1 \mreg/_08015_ ( .A(\mreg/_04534_ ), .ZN(\mreg/_02121_ ) );
OAI21_X1 \mreg/_08016_ ( .A(\mreg/_02120_ ), .B1(\mreg/_01678_ ), .B2(\mreg/_02121_ ), .ZN(\mreg/_02122_ ) );
AOI221_X4 \mreg/_08017_ ( .A(\mreg/_02122_ ), .B1(\mreg/_04470_ ), .B2(\mreg/_01195_ ), .C1(\mreg/_04438_ ), .C2(\mreg/_01660_ ), .ZN(\mreg/_02123_ ) );
NAND3_X1 \mreg/_08018_ ( .A1(\mreg/_01398_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04374_ ), .ZN(\mreg/_02124_ ) );
NAND3_X1 \mreg/_08019_ ( .A1(\mreg/_01496_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04406_ ), .ZN(\mreg/_02125_ ) );
NAND2_X1 \mreg/_08020_ ( .A1(\mreg/_02124_ ), .A2(\mreg/_02125_ ), .ZN(\mreg/_02126_ ) );
AOI221_X4 \mreg/_08021_ ( .A(\mreg/_02126_ ), .B1(\mreg/_04342_ ), .B2(\mreg/_01611_ ), .C1(\mreg/_04310_ ), .C2(\mreg/_01499_ ), .ZN(\mreg/_02127_ ) );
NAND3_X1 \mreg/_08022_ ( .A1(\mreg/_01082_ ), .A2(\mreg/_04150_ ), .A3(\mreg/_01981_ ), .ZN(\mreg/_02128_ ) );
NAND3_X1 \mreg/_08023_ ( .A1(\mreg/_01621_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04182_ ), .ZN(\mreg/_02129_ ) );
NAND4_X1 \mreg/_08024_ ( .A1(\mreg/_01667_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04214_ ), .A4(\mreg/_01212_ ), .ZN(\mreg/_02130_ ) );
NAND4_X1 \mreg/_08025_ ( .A1(\mreg/_01211_ ), .A2(\mreg/_01981_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04246_ ), .ZN(\mreg/_02131_ ) );
AND4_X1 \mreg/_08026_ ( .A1(\mreg/_02128_ ), .A2(\mreg/_02129_ ), .A3(\mreg/_02130_ ), .A4(\mreg/_02131_ ), .ZN(\mreg/_02132_ ) );
AND4_X4 \mreg/_08027_ ( .A1(\mreg/_02119_ ), .A2(\mreg/_02123_ ), .A3(\mreg/_02127_ ), .A4(\mreg/_02132_ ), .ZN(\mreg/_02133_ ) );
NAND3_X1 \mreg/_08028_ ( .A1(\mreg/_01059_ ), .A2(\mreg/_01277_ ), .A3(\mreg/_04790_ ), .ZN(\mreg/_02134_ ) );
AND3_X1 \mreg/_08029_ ( .A1(\mreg/_01072_ ), .A2(\mreg/_01357_ ), .A3(\mreg/_04278_ ), .ZN(\mreg/_02135_ ) );
AOI221_X4 \mreg/_08030_ ( .A(\mreg/_02135_ ), .B1(\mreg/_01105_ ), .B2(\mreg/_04726_ ), .C1(\mreg/_04630_ ), .C2(\mreg/_01221_ ), .ZN(\mreg/_02136_ ) );
NAND3_X1 \mreg/_08031_ ( .A1(\mreg/_01292_ ), .A2(\mreg/_01087_ ), .A3(\mreg/_04758_ ), .ZN(\mreg/_02137_ ) );
AND3_X1 \mreg/_08032_ ( .A1(\mreg/_01380_ ), .A2(\mreg/_01133_ ), .A3(\mreg/_04854_ ), .ZN(\mreg/_02138_ ) );
AOI21_X1 \mreg/_08033_ ( .A(\mreg/_02138_ ), .B1(\mreg/_04822_ ), .B2(\mreg/_01431_ ), .ZN(\mreg/_02139_ ) );
AND4_X1 \mreg/_08034_ ( .A1(\mreg/_02134_ ), .A2(\mreg/_02136_ ), .A3(\mreg/_02137_ ), .A4(\mreg/_02139_ ), .ZN(\mreg/_02140_ ) );
NAND3_X1 \mreg/_08035_ ( .A1(\mreg/_01155_ ), .A2(\mreg/_01436_ ), .A3(\mreg/_04918_ ), .ZN(\mreg/_02141_ ) );
NAND3_X1 \mreg/_08036_ ( .A1(\mreg/_01159_ ), .A2(\mreg/_01282_ ), .A3(\mreg/_03958_ ), .ZN(\mreg/_02142_ ) );
NAND3_X1 \mreg/_08037_ ( .A1(\mreg/_01292_ ), .A2(\mreg/_01293_ ), .A3(\mreg/_04886_ ), .ZN(\mreg/_02143_ ) );
NAND3_X1 \mreg/_08038_ ( .A1(\mreg/_01165_ ), .A2(\mreg/_01477_ ), .A3(\mreg/_03990_ ), .ZN(\mreg/_02144_ ) );
AND4_X1 \mreg/_08039_ ( .A1(\mreg/_02141_ ), .A2(\mreg/_02142_ ), .A3(\mreg/_02143_ ), .A4(\mreg/_02144_ ), .ZN(\mreg/_02145_ ) );
NAND3_X1 \mreg/_08040_ ( .A1(\mreg/_01298_ ), .A2(\mreg/_04022_ ), .A3(\mreg/_01299_ ), .ZN(\mreg/_02146_ ) );
NAND3_X1 \mreg/_08041_ ( .A1(\mreg/_01301_ ), .A2(\mreg/_01302_ ), .A3(\mreg/_04086_ ), .ZN(\mreg/_02147_ ) );
NAND3_X1 \mreg/_08042_ ( .A1(\mreg/_01235_ ), .A2(\mreg/_01295_ ), .A3(\mreg/_04054_ ), .ZN(\mreg/_02148_ ) );
NAND3_X1 \mreg/_08043_ ( .A1(\mreg/_01308_ ), .A2(\mreg/_01309_ ), .A3(\mreg/_04118_ ), .ZN(\mreg/_02149_ ) );
AND4_X1 \mreg/_08044_ ( .A1(\mreg/_02146_ ), .A2(\mreg/_02147_ ), .A3(\mreg/_02148_ ), .A4(\mreg/_02149_ ), .ZN(\mreg/_02150_ ) );
NAND4_X1 \mreg/_08045_ ( .A1(\mreg/_02133_ ), .A2(\mreg/_02140_ ), .A3(\mreg/_02145_ ), .A4(\mreg/_02150_ ), .ZN(\mreg/_03926_ ) );
NAND3_X1 \mreg/_08046_ ( .A1(\mreg/_01083_ ), .A2(\mreg/_04567_ ), .A3(\mreg/_01597_ ), .ZN(\mreg/_02151_ ) );
NAND3_X1 \mreg/_08047_ ( .A1(\mreg/_01143_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04663_ ), .ZN(\mreg/_02152_ ) );
NAND3_X1 \mreg/_08048_ ( .A1(\mreg/_01148_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04599_ ), .ZN(\mreg/_02153_ ) );
INV_X1 \mreg/_08049_ ( .A(\mreg/_00055_ ), .ZN(\mreg/_02154_ ) );
NAND3_X1 \mreg/_08050_ ( .A1(\mreg/_01140_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_02154_ ), .ZN(\mreg/_02155_ ) );
AND4_X1 \mreg/_08051_ ( .A1(\mreg/_02151_ ), .A2(\mreg/_02152_ ), .A3(\mreg/_02153_ ), .A4(\mreg/_02155_ ), .ZN(\mreg/_02156_ ) );
NAND3_X1 \mreg/_08052_ ( .A1(\mreg/_01091_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04375_ ), .ZN(\mreg/_02157_ ) );
NAND3_X1 \mreg/_08053_ ( .A1(\mreg/_01097_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04407_ ), .ZN(\mreg/_02158_ ) );
NAND2_X1 \mreg/_08054_ ( .A1(\mreg/_02157_ ), .A2(\mreg/_02158_ ), .ZN(\mreg/_02159_ ) );
AOI221_X4 \mreg/_08055_ ( .A(\mreg/_02159_ ), .B1(\mreg/_04343_ ), .B2(\mreg/_01205_ ), .C1(\mreg/_04311_ ), .C2(\mreg/_01207_ ), .ZN(\mreg/_02160_ ) );
NAND3_X1 \mreg/_08056_ ( .A1(\mreg/_01121_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04471_ ), .ZN(\mreg/_02161_ ) );
NAND3_X1 \mreg/_08057_ ( .A1(\mreg/_01082_ ), .A2(\mreg/_04439_ ), .A3(\mreg/_01162_ ), .ZN(\mreg/_02162_ ) );
NAND4_X1 \mreg/_08058_ ( .A1(\mreg/_01667_ ), .A2(\mreg/_01162_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04503_ ), .ZN(\mreg/_02163_ ) );
NAND4_X1 \mreg/_08059_ ( .A1(\mreg/_01162_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_01211_ ), .A4(\mreg/_04535_ ), .ZN(\mreg/_02164_ ) );
AND4_X1 \mreg/_08060_ ( .A1(\mreg/_02161_ ), .A2(\mreg/_02162_ ), .A3(\mreg/_02163_ ), .A4(\mreg/_02164_ ), .ZN(\mreg/_02165_ ) );
NAND4_X1 \mreg/_08061_ ( .A1(\mreg/_01501_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04215_ ), .A4(\mreg/_01372_ ), .ZN(\mreg/_02166_ ) );
INV_X1 \mreg/_08062_ ( .A(\mreg/_04247_ ), .ZN(\mreg/_02167_ ) );
OAI21_X1 \mreg/_08063_ ( .A(\mreg/_02166_ ), .B1(\mreg/_01374_ ), .B2(\mreg/_02167_ ), .ZN(\mreg/_02168_ ) );
AOI221_X4 \mreg/_08064_ ( .A(\mreg/_02168_ ), .B1(\mreg/_04183_ ), .B2(\mreg/_01465_ ), .C1(\mreg/_04151_ ), .C2(\mreg/_01505_ ), .ZN(\mreg/_02169_ ) );
AND4_X2 \mreg/_08065_ ( .A1(\mreg/_02156_ ), .A2(\mreg/_02160_ ), .A3(\mreg/_02165_ ), .A4(\mreg/_02169_ ), .ZN(\mreg/_02170_ ) );
NAND3_X1 \mreg/_08066_ ( .A1(\mreg/_01059_ ), .A2(\mreg/_01287_ ), .A3(\mreg/_04791_ ), .ZN(\mreg/_02171_ ) );
AND3_X1 \mreg/_08067_ ( .A1(\mreg/_01072_ ), .A2(\mreg/_01357_ ), .A3(\mreg/_04279_ ), .ZN(\mreg/_02172_ ) );
AOI221_X4 \mreg/_08068_ ( .A(\mreg/_02172_ ), .B1(\mreg/_01105_ ), .B2(\mreg/_04727_ ), .C1(\mreg/_04631_ ), .C2(\mreg/_01221_ ), .ZN(\mreg/_02173_ ) );
NAND3_X1 \mreg/_08069_ ( .A1(\mreg/_01292_ ), .A2(\mreg/_01087_ ), .A3(\mreg/_04759_ ), .ZN(\mreg/_02174_ ) );
AND3_X1 \mreg/_08070_ ( .A1(\mreg/_01380_ ), .A2(\mreg/_01133_ ), .A3(\mreg/_04855_ ), .ZN(\mreg/_02175_ ) );
AOI21_X1 \mreg/_08071_ ( .A(\mreg/_02175_ ), .B1(\mreg/_04823_ ), .B2(\mreg/_01431_ ), .ZN(\mreg/_02176_ ) );
AND4_X1 \mreg/_08072_ ( .A1(\mreg/_02171_ ), .A2(\mreg/_02173_ ), .A3(\mreg/_02174_ ), .A4(\mreg/_02176_ ), .ZN(\mreg/_02177_ ) );
NAND3_X1 \mreg/_08073_ ( .A1(\mreg/_01155_ ), .A2(\mreg/_01436_ ), .A3(\mreg/_04919_ ), .ZN(\mreg/_02178_ ) );
NAND3_X1 \mreg/_08074_ ( .A1(\mreg/_01159_ ), .A2(\mreg/_01282_ ), .A3(\mreg/_03959_ ), .ZN(\mreg/_02179_ ) );
NAND3_X1 \mreg/_08075_ ( .A1(\mreg/_01339_ ), .A2(\mreg/_01293_ ), .A3(\mreg/_04887_ ), .ZN(\mreg/_02180_ ) );
NAND3_X1 \mreg/_08076_ ( .A1(\mreg/_01165_ ), .A2(\mreg/_01477_ ), .A3(\mreg/_03991_ ), .ZN(\mreg/_02181_ ) );
AND4_X1 \mreg/_08077_ ( .A1(\mreg/_02178_ ), .A2(\mreg/_02179_ ), .A3(\mreg/_02180_ ), .A4(\mreg/_02181_ ), .ZN(\mreg/_02182_ ) );
NAND3_X1 \mreg/_08078_ ( .A1(\mreg/_01298_ ), .A2(\mreg/_04023_ ), .A3(\mreg/_01242_ ), .ZN(\mreg/_02183_ ) );
NAND3_X1 \mreg/_08079_ ( .A1(\mreg/_01301_ ), .A2(\mreg/_01306_ ), .A3(\mreg/_04087_ ), .ZN(\mreg/_02184_ ) );
NAND3_X1 \mreg/_08080_ ( .A1(\mreg/_01235_ ), .A2(\mreg/_01295_ ), .A3(\mreg/_04055_ ), .ZN(\mreg/_02185_ ) );
NAND3_X1 \mreg/_08081_ ( .A1(\mreg/_01308_ ), .A2(\mreg/_01309_ ), .A3(\mreg/_04119_ ), .ZN(\mreg/_02186_ ) );
AND4_X1 \mreg/_08082_ ( .A1(\mreg/_02183_ ), .A2(\mreg/_02184_ ), .A3(\mreg/_02185_ ), .A4(\mreg/_02186_ ), .ZN(\mreg/_02187_ ) );
NAND4_X1 \mreg/_08083_ ( .A1(\mreg/_02170_ ), .A2(\mreg/_02177_ ), .A3(\mreg/_02182_ ), .A4(\mreg/_02187_ ), .ZN(\mreg/_03927_ ) );
NAND3_X1 \mreg/_08084_ ( .A1(\mreg/_01125_ ), .A2(\mreg/_01086_ ), .A3(\mreg/_04760_ ), .ZN(\mreg/_02188_ ) );
INV_X1 \mreg/_08085_ ( .A(\mreg/_04728_ ), .ZN(\mreg/_02189_ ) );
OAI21_X1 \mreg/_08086_ ( .A(\mreg/_02188_ ), .B1(\mreg/_01786_ ), .B2(\mreg/_02189_ ), .ZN(\mreg/_02190_ ) );
AOI221_X4 \mreg/_08087_ ( .A(\mreg/_02190_ ), .B1(\mreg/_04824_ ), .B2(\mreg/_01430_ ), .C1(\mreg/_04792_ ), .C2(\mreg/_01228_ ), .ZN(\mreg/_02191_ ) );
NAND3_X1 \mreg/_08088_ ( .A1(\mreg/_01139_ ), .A2(\mreg/_01108_ ), .A3(\mreg/_04120_ ), .ZN(\mreg/_02192_ ) );
INV_X1 \mreg/_08089_ ( .A(\mreg/_04056_ ), .ZN(\mreg/_02193_ ) );
OAI21_X1 \mreg/_08090_ ( .A(\mreg/_02192_ ), .B1(\mreg/_01791_ ), .B2(\mreg/_02193_ ), .ZN(\mreg/_02194_ ) );
AOI221_X1 \mreg/_08091_ ( .A(\mreg/_02194_ ), .B1(\mreg/_03960_ ), .B2(\mreg/_01361_ ), .C1(\mreg/_04920_ ), .C2(\mreg/_01362_ ), .ZN(\mreg/_02195_ ) );
NAND4_X1 \mreg/_08092_ ( .A1(\mreg/_01365_ ), .A2(\mreg/_01116_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04504_ ), .ZN(\mreg/_02196_ ) );
INV_X1 \mreg/_08093_ ( .A(\mreg/_04536_ ), .ZN(\mreg/_02197_ ) );
OAI21_X1 \mreg/_08094_ ( .A(\mreg/_02196_ ), .B1(\mreg/_01190_ ), .B2(\mreg/_02197_ ), .ZN(\mreg/_02198_ ) );
INV_X1 \mreg/_08095_ ( .A(\mreg/_00056_ ), .ZN(\mreg/_02199_ ) );
AOI221_X1 \mreg/_08096_ ( .A(\mreg/_02198_ ), .B1(\mreg/_02199_ ), .B2(\mreg/_01172_ ), .C1(\mreg/_04664_ ), .C2(\mreg/_01174_ ), .ZN(\mreg/_02200_ ) );
NAND4_X1 \mreg/_08097_ ( .A1(\mreg/_01089_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04216_ ), .A4(\mreg/_01062_ ), .ZN(\mreg/_02201_ ) );
INV_X1 \mreg/_08098_ ( .A(\mreg/_04248_ ), .ZN(\mreg/_02202_ ) );
OAI21_X1 \mreg/_08099_ ( .A(\mreg/_02201_ ), .B1(\mreg/_01068_ ), .B2(\mreg/_02202_ ), .ZN(\mreg/_02203_ ) );
AOI221_X4 \mreg/_08100_ ( .A(\mreg/_02203_ ), .B1(\mreg/_04344_ ), .B2(\mreg/_01204_ ), .C1(\mreg/_04312_ ), .C2(\mreg/_01206_ ), .ZN(\mreg/_02204_ ) );
NAND4_X1 \mreg/_08101_ ( .A1(\mreg/_02191_ ), .A2(\mreg/_02195_ ), .A3(\mreg/_02200_ ), .A4(\mreg/_02204_ ), .ZN(\mreg/_02205_ ) );
NAND3_X1 \mreg/_08102_ ( .A1(\mreg/_01381_ ), .A2(\mreg/_01239_ ), .A3(\mreg/_04856_ ), .ZN(\mreg/_02206_ ) );
NAND3_X1 \mreg/_08103_ ( .A1(\mreg/_01621_ ), .A2(\mreg/_01387_ ), .A3(\mreg/_04280_ ), .ZN(\mreg/_02207_ ) );
NAND3_X1 \mreg/_08104_ ( .A1(\mreg/_01386_ ), .A2(\mreg/_01248_ ), .A3(\mreg/_04632_ ), .ZN(\mreg/_02208_ ) );
NAND3_X1 \mreg/_08105_ ( .A1(\mreg/_01250_ ), .A2(\mreg/_01251_ ), .A3(\mreg/_04888_ ), .ZN(\mreg/_02209_ ) );
NAND4_X1 \mreg/_08106_ ( .A1(\mreg/_02206_ ), .A2(\mreg/_02207_ ), .A3(\mreg/_02208_ ), .A4(\mreg/_02209_ ), .ZN(\mreg/_02210_ ) );
NAND3_X1 \mreg/_08107_ ( .A1(\mreg/_01291_ ), .A2(\mreg/_04024_ ), .A3(\mreg/_01391_ ), .ZN(\mreg/_02211_ ) );
INV_X1 \mreg/_08108_ ( .A(\mreg/_04088_ ), .ZN(\mreg/_02212_ ) );
INV_X1 \mreg/_08109_ ( .A(\mreg/_03992_ ), .ZN(\mreg/_02213_ ) );
OAI221_X1 \mreg/_08110_ ( .A(\mreg/_02211_ ), .B1(\mreg/_01393_ ), .B2(\mreg/_02212_ ), .C1(\mreg/_02213_ ), .C2(\mreg/_01396_ ), .ZN(\mreg/_02214_ ) );
NAND3_X2 \mreg/_08111_ ( .A1(\mreg/_01398_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04376_ ), .ZN(\mreg/_02215_ ) );
NAND3_X2 \mreg/_08112_ ( .A1(\mreg/_01096_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04408_ ), .ZN(\mreg/_02216_ ) );
NAND2_X1 \mreg/_08113_ ( .A1(\mreg/_02215_ ), .A2(\mreg/_02216_ ), .ZN(\mreg/_02217_ ) );
AOI221_X2 \mreg/_08114_ ( .A(\mreg/_02217_ ), .B1(\mreg/_04184_ ), .B2(\mreg/_01074_ ), .C1(\mreg/_04152_ ), .C2(\mreg/_01079_ ), .ZN(\mreg/_02218_ ) );
AND3_X1 \mreg/_08115_ ( .A1(\mreg/_01255_ ), .A2(\mreg/_04440_ ), .A3(\mreg/_01127_ ), .ZN(\mreg/_02219_ ) );
AOI21_X1 \mreg/_08116_ ( .A(\mreg/_02219_ ), .B1(\mreg/_01196_ ), .B2(\mreg/_04472_ ), .ZN(\mreg/_02220_ ) );
NAND3_X1 \mreg/_08117_ ( .A1(\mreg/_01177_ ), .A2(\mreg/_04568_ ), .A3(\mreg/_01178_ ), .ZN(\mreg/_02221_ ) );
NAND3_X1 \mreg/_08118_ ( .A1(\mreg/_01304_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04600_ ), .ZN(\mreg/_02222_ ) );
NAND4_X4 \mreg/_08119_ ( .A1(\mreg/_02218_ ), .A2(\mreg/_02220_ ), .A3(\mreg/_02221_ ), .A4(\mreg/_02222_ ), .ZN(\mreg/_02223_ ) );
OR4_X2 \mreg/_08120_ ( .A1(\mreg/_02205_ ), .A2(\mreg/_02210_ ), .A3(\mreg/_02214_ ), .A4(\mreg/_02223_ ), .ZN(\mreg/_03928_ ) );
NAND3_X1 \mreg/_08121_ ( .A1(\mreg/_01083_ ), .A2(\mreg/_04569_ ), .A3(\mreg/_01597_ ), .ZN(\mreg/_02224_ ) );
NAND3_X1 \mreg/_08122_ ( .A1(\mreg/_01143_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04665_ ), .ZN(\mreg/_02225_ ) );
NAND3_X1 \mreg/_08123_ ( .A1(\mreg/_01148_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04601_ ), .ZN(\mreg/_02226_ ) );
INV_X1 \mreg/_08124_ ( .A(\mreg/_00057_ ), .ZN(\mreg/_02227_ ) );
NAND3_X1 \mreg/_08125_ ( .A1(\mreg/_01140_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_02227_ ), .ZN(\mreg/_02228_ ) );
AND4_X1 \mreg/_08126_ ( .A1(\mreg/_02224_ ), .A2(\mreg/_02225_ ), .A3(\mreg/_02226_ ), .A4(\mreg/_02228_ ), .ZN(\mreg/_02229_ ) );
NAND4_X1 \mreg/_08127_ ( .A1(\mreg/_01269_ ), .A2(\mreg/_01366_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04505_ ), .ZN(\mreg/_02230_ ) );
INV_X1 \mreg/_08128_ ( .A(\mreg/_04537_ ), .ZN(\mreg/_02231_ ) );
OAI21_X1 \mreg/_08129_ ( .A(\mreg/_02230_ ), .B1(\mreg/_01678_ ), .B2(\mreg/_02231_ ), .ZN(\mreg/_02232_ ) );
AOI221_X1 \mreg/_08130_ ( .A(\mreg/_02232_ ), .B1(\mreg/_04473_ ), .B2(\mreg/_01195_ ), .C1(\mreg/_04441_ ), .C2(\mreg/_01660_ ), .ZN(\mreg/_02233_ ) );
NAND3_X1 \mreg/_08131_ ( .A1(\mreg/_01398_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04377_ ), .ZN(\mreg/_02234_ ) );
NAND3_X1 \mreg/_08132_ ( .A1(\mreg/_01096_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04409_ ), .ZN(\mreg/_02235_ ) );
NAND2_X1 \mreg/_08133_ ( .A1(\mreg/_02234_ ), .A2(\mreg/_02235_ ), .ZN(\mreg/_02236_ ) );
AOI221_X4 \mreg/_08134_ ( .A(\mreg/_02236_ ), .B1(\mreg/_04345_ ), .B2(\mreg/_01611_ ), .C1(\mreg/_04313_ ), .C2(\mreg/_01377_ ), .ZN(\mreg/_02237_ ) );
NAND3_X1 \mreg/_08135_ ( .A1(\mreg/_01082_ ), .A2(\mreg/_04153_ ), .A3(\mreg/_01981_ ), .ZN(\mreg/_02238_ ) );
NAND3_X1 \mreg/_08136_ ( .A1(\mreg/_01621_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04185_ ), .ZN(\mreg/_02239_ ) );
NAND4_X1 \mreg/_08137_ ( .A1(\mreg/_01667_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04217_ ), .A4(\mreg/_01212_ ), .ZN(\mreg/_02240_ ) );
NAND4_X1 \mreg/_08138_ ( .A1(\mreg/_01211_ ), .A2(\mreg/_01981_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04249_ ), .ZN(\mreg/_02241_ ) );
AND4_X1 \mreg/_08139_ ( .A1(\mreg/_02238_ ), .A2(\mreg/_02239_ ), .A3(\mreg/_02240_ ), .A4(\mreg/_02241_ ), .ZN(\mreg/_02242_ ) );
AND4_X1 \mreg/_08140_ ( .A1(\mreg/_02229_ ), .A2(\mreg/_02233_ ), .A3(\mreg/_02237_ ), .A4(\mreg/_02242_ ), .ZN(\mreg/_02243_ ) );
NAND3_X1 \mreg/_08141_ ( .A1(\mreg/_01059_ ), .A2(\mreg/_01287_ ), .A3(\mreg/_04793_ ), .ZN(\mreg/_02244_ ) );
AND3_X1 \mreg/_08142_ ( .A1(\mreg/_01072_ ), .A2(\mreg/_01357_ ), .A3(\mreg/_04281_ ), .ZN(\mreg/_02245_ ) );
AOI221_X4 \mreg/_08143_ ( .A(\mreg/_02245_ ), .B1(\mreg/_01105_ ), .B2(\mreg/_04729_ ), .C1(\mreg/_04633_ ), .C2(\mreg/_01221_ ), .ZN(\mreg/_02246_ ) );
NAND3_X1 \mreg/_08144_ ( .A1(\mreg/_01292_ ), .A2(\mreg/_01087_ ), .A3(\mreg/_04761_ ), .ZN(\mreg/_02247_ ) );
AND3_X1 \mreg/_08145_ ( .A1(\mreg/_01380_ ), .A2(\mreg/_01133_ ), .A3(\mreg/_04857_ ), .ZN(\mreg/_02248_ ) );
AOI21_X1 \mreg/_08146_ ( .A(\mreg/_02248_ ), .B1(\mreg/_04825_ ), .B2(\mreg/_01431_ ), .ZN(\mreg/_02249_ ) );
AND4_X1 \mreg/_08147_ ( .A1(\mreg/_02244_ ), .A2(\mreg/_02246_ ), .A3(\mreg/_02247_ ), .A4(\mreg/_02249_ ), .ZN(\mreg/_02250_ ) );
NAND3_X1 \mreg/_08148_ ( .A1(\mreg/_01155_ ), .A2(\mreg/_01436_ ), .A3(\mreg/_04921_ ), .ZN(\mreg/_02251_ ) );
NAND3_X1 \mreg/_08149_ ( .A1(\mreg/_01158_ ), .A2(\mreg/_01282_ ), .A3(\mreg/_03961_ ), .ZN(\mreg/_02252_ ) );
NAND3_X1 \mreg/_08150_ ( .A1(\mreg/_01339_ ), .A2(\mreg/_01293_ ), .A3(\mreg/_04889_ ), .ZN(\mreg/_02253_ ) );
NAND3_X1 \mreg/_08151_ ( .A1(\mreg/_01113_ ), .A2(\mreg/_01477_ ), .A3(\mreg/_03993_ ), .ZN(\mreg/_02254_ ) );
AND4_X1 \mreg/_08152_ ( .A1(\mreg/_02251_ ), .A2(\mreg/_02252_ ), .A3(\mreg/_02253_ ), .A4(\mreg/_02254_ ), .ZN(\mreg/_02255_ ) );
NAND3_X1 \mreg/_08153_ ( .A1(\mreg/_01298_ ), .A2(\mreg/_04025_ ), .A3(\mreg/_01242_ ), .ZN(\mreg/_02256_ ) );
NAND3_X1 \mreg/_08154_ ( .A1(\mreg/_01301_ ), .A2(\mreg/_01306_ ), .A3(\mreg/_04089_ ), .ZN(\mreg/_02257_ ) );
NAND3_X1 \mreg/_08155_ ( .A1(\mreg/_01235_ ), .A2(\mreg/_01295_ ), .A3(\mreg/_04057_ ), .ZN(\mreg/_02258_ ) );
NAND3_X1 \mreg/_08156_ ( .A1(\mreg/_01308_ ), .A2(\mreg/_01309_ ), .A3(\mreg/_04121_ ), .ZN(\mreg/_02259_ ) );
AND4_X1 \mreg/_08157_ ( .A1(\mreg/_02256_ ), .A2(\mreg/_02257_ ), .A3(\mreg/_02258_ ), .A4(\mreg/_02259_ ), .ZN(\mreg/_02260_ ) );
NAND4_X1 \mreg/_08158_ ( .A1(\mreg/_02243_ ), .A2(\mreg/_02250_ ), .A3(\mreg/_02255_ ), .A4(\mreg/_02260_ ), .ZN(\mreg/_03929_ ) );
NAND3_X1 \mreg/_08159_ ( .A1(\mreg/_01083_ ), .A2(\mreg/_04570_ ), .A3(\mreg/_01597_ ), .ZN(\mreg/_02261_ ) );
NAND3_X1 \mreg/_08160_ ( .A1(\mreg/_01143_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04666_ ), .ZN(\mreg/_02262_ ) );
NAND3_X1 \mreg/_08161_ ( .A1(\mreg/_01148_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04602_ ), .ZN(\mreg/_02263_ ) );
INV_X1 \mreg/_08162_ ( .A(\mreg/_00058_ ), .ZN(\mreg/_02264_ ) );
NAND3_X1 \mreg/_08163_ ( .A1(\mreg/_01140_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_02264_ ), .ZN(\mreg/_02265_ ) );
AND4_X1 \mreg/_08164_ ( .A1(\mreg/_02261_ ), .A2(\mreg/_02262_ ), .A3(\mreg/_02263_ ), .A4(\mreg/_02265_ ), .ZN(\mreg/_02266_ ) );
NAND4_X1 \mreg/_08165_ ( .A1(\mreg/_01269_ ), .A2(\mreg/_01366_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04506_ ), .ZN(\mreg/_02267_ ) );
INV_X1 \mreg/_08166_ ( .A(\mreg/_04538_ ), .ZN(\mreg/_02268_ ) );
OAI21_X1 \mreg/_08167_ ( .A(\mreg/_02267_ ), .B1(\mreg/_01678_ ), .B2(\mreg/_02268_ ), .ZN(\mreg/_02269_ ) );
AOI221_X4 \mreg/_08168_ ( .A(\mreg/_02269_ ), .B1(\mreg/_04474_ ), .B2(\mreg/_01195_ ), .C1(\mreg/_04442_ ), .C2(\mreg/_01660_ ), .ZN(\mreg/_02270_ ) );
NAND3_X1 \mreg/_08169_ ( .A1(\mreg/_01398_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04378_ ), .ZN(\mreg/_02271_ ) );
NAND3_X1 \mreg/_08170_ ( .A1(\mreg/_01096_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04410_ ), .ZN(\mreg/_02272_ ) );
NAND2_X1 \mreg/_08171_ ( .A1(\mreg/_02271_ ), .A2(\mreg/_02272_ ), .ZN(\mreg/_02273_ ) );
AOI221_X4 \mreg/_08172_ ( .A(\mreg/_02273_ ), .B1(\mreg/_04346_ ), .B2(\mreg/_01204_ ), .C1(\mreg/_04314_ ), .C2(\mreg/_01377_ ), .ZN(\mreg/_02274_ ) );
NAND4_X1 \mreg/_08173_ ( .A1(\mreg/_01501_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04218_ ), .A4(\mreg/_01372_ ), .ZN(\mreg/_02275_ ) );
INV_X1 \mreg/_08174_ ( .A(\mreg/_04250_ ), .ZN(\mreg/_02276_ ) );
OAI21_X1 \mreg/_08175_ ( .A(\mreg/_02275_ ), .B1(\mreg/_01374_ ), .B2(\mreg/_02276_ ), .ZN(\mreg/_02277_ ) );
AOI221_X4 \mreg/_08176_ ( .A(\mreg/_02277_ ), .B1(\mreg/_04186_ ), .B2(\mreg/_01465_ ), .C1(\mreg/_04154_ ), .C2(\mreg/_01505_ ), .ZN(\mreg/_02278_ ) );
AND4_X2 \mreg/_08177_ ( .A1(\mreg/_02266_ ), .A2(\mreg/_02270_ ), .A3(\mreg/_02274_ ), .A4(\mreg/_02278_ ), .ZN(\mreg/_02279_ ) );
NAND3_X1 \mreg/_08178_ ( .A1(\mreg/_01383_ ), .A2(\mreg/_01287_ ), .A3(\mreg/_04282_ ), .ZN(\mreg/_02280_ ) );
AND3_X1 \mreg/_08179_ ( .A1(\mreg/_01098_ ), .A2(\mreg/_01144_ ), .A3(\mreg/_04858_ ), .ZN(\mreg/_02281_ ) );
AOI21_X1 \mreg/_08180_ ( .A(\mreg/_02281_ ), .B1(\mreg/_04826_ ), .B2(\mreg/_01431_ ), .ZN(\mreg/_02282_ ) );
AOI22_X1 \mreg/_08181_ ( .A1(\mreg/_04634_ ), .A2(\mreg/_01222_ ), .B1(\mreg/_01219_ ), .B2(\mreg/_04730_ ), .ZN(\mreg/_02283_ ) );
AOI22_X1 \mreg/_08182_ ( .A1(\mreg/_01284_ ), .A2(\mreg/_04794_ ), .B1(\mreg/_04762_ ), .B2(\mreg/_01229_ ), .ZN(\mreg/_02284_ ) );
AND4_X1 \mreg/_08183_ ( .A1(\mreg/_02280_ ), .A2(\mreg/_02282_ ), .A3(\mreg/_02283_ ), .A4(\mreg/_02284_ ), .ZN(\mreg/_02285_ ) );
AND3_X1 \mreg/_08184_ ( .A1(\mreg/_01113_ ), .A2(\mreg/_01309_ ), .A3(\mreg/_03994_ ), .ZN(\mreg/_02286_ ) );
AND3_X1 \mreg/_08185_ ( .A1(\mreg/_01158_ ), .A2(\mreg/_01239_ ), .A3(\mreg/_03962_ ), .ZN(\mreg/_02287_ ) );
AND3_X1 \mreg/_08186_ ( .A1(\mreg/_01155_ ), .A2(\mreg/_01387_ ), .A3(\mreg/_04922_ ), .ZN(\mreg/_02288_ ) );
AND3_X1 \mreg/_08187_ ( .A1(\mreg/_01250_ ), .A2(\mreg/_04890_ ), .A3(\mreg/_01251_ ), .ZN(\mreg/_02289_ ) );
NOR4_X1 \mreg/_08188_ ( .A1(\mreg/_02286_ ), .A2(\mreg/_02287_ ), .A3(\mreg/_02288_ ), .A4(\mreg/_02289_ ), .ZN(\mreg/_02290_ ) );
NAND3_X1 \mreg/_08189_ ( .A1(\mreg/_01298_ ), .A2(\mreg/_04026_ ), .A3(\mreg/_01242_ ), .ZN(\mreg/_02291_ ) );
NAND3_X1 \mreg/_08190_ ( .A1(\mreg/_01232_ ), .A2(\mreg/_01306_ ), .A3(\mreg/_04090_ ), .ZN(\mreg/_02292_ ) );
NAND3_X1 \mreg/_08191_ ( .A1(\mreg/_01235_ ), .A2(\mreg/_01295_ ), .A3(\mreg/_04058_ ), .ZN(\mreg/_02293_ ) );
NAND3_X1 \mreg/_08192_ ( .A1(\mreg/_01238_ ), .A2(\mreg/_01309_ ), .A3(\mreg/_04122_ ), .ZN(\mreg/_02294_ ) );
AND4_X1 \mreg/_08193_ ( .A1(\mreg/_02291_ ), .A2(\mreg/_02292_ ), .A3(\mreg/_02293_ ), .A4(\mreg/_02294_ ), .ZN(\mreg/_02295_ ) );
NAND4_X1 \mreg/_08194_ ( .A1(\mreg/_02279_ ), .A2(\mreg/_02285_ ), .A3(\mreg/_02290_ ), .A4(\mreg/_02295_ ), .ZN(\mreg/_03930_ ) );
NAND3_X1 \mreg/_08195_ ( .A1(\mreg/_01147_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04603_ ), .ZN(\mreg/_02296_ ) );
NAND3_X1 \mreg/_08196_ ( .A1(\mreg/_01255_ ), .A2(\mreg/_04571_ ), .A3(\mreg/_01150_ ), .ZN(\mreg/_02297_ ) );
NAND2_X1 \mreg/_08197_ ( .A1(\mreg/_02296_ ), .A2(\mreg/_02297_ ), .ZN(\mreg/_02298_ ) );
INV_X1 \mreg/_08198_ ( .A(\mreg/_00059_ ), .ZN(\mreg/_02299_ ) );
AOI221_X4 \mreg/_08199_ ( .A(\mreg/_02298_ ), .B1(\mreg/_02299_ ), .B2(\mreg/_01172_ ), .C1(\mreg/_04667_ ), .C2(\mreg/_01175_ ), .ZN(\mreg/_02300_ ) );
NAND3_X1 \mreg/_08200_ ( .A1(\mreg/_01091_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04379_ ), .ZN(\mreg/_02301_ ) );
NAND3_X1 \mreg/_08201_ ( .A1(\mreg/_01097_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04411_ ), .ZN(\mreg/_02302_ ) );
NAND2_X1 \mreg/_08202_ ( .A1(\mreg/_02301_ ), .A2(\mreg/_02302_ ), .ZN(\mreg/_02303_ ) );
AOI221_X4 \mreg/_08203_ ( .A(\mreg/_02303_ ), .B1(\mreg/_04347_ ), .B2(\mreg/_01205_ ), .C1(\mreg/_04315_ ), .C2(\mreg/_01207_ ), .ZN(\mreg/_02304_ ) );
NAND4_X1 \mreg/_08204_ ( .A1(\mreg/_01188_ ), .A2(\mreg/_01161_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04507_ ), .ZN(\mreg/_02305_ ) );
NAND4_X1 \mreg/_08205_ ( .A1(\mreg/_01161_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_01211_ ), .A4(\mreg/_04539_ ), .ZN(\mreg/_02306_ ) );
NAND2_X1 \mreg/_08206_ ( .A1(\mreg/_02305_ ), .A2(\mreg/_02306_ ), .ZN(\mreg/_02307_ ) );
AOI221_X4 \mreg/_08207_ ( .A(\mreg/_02307_ ), .B1(\mreg/_01660_ ), .B2(\mreg/_04443_ ), .C1(\mreg/_04475_ ), .C2(\mreg/_01196_ ), .ZN(\mreg/_02308_ ) );
NAND4_X1 \mreg/_08208_ ( .A1(\mreg/_01501_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04219_ ), .A4(\mreg/_01372_ ), .ZN(\mreg/_02309_ ) );
INV_X1 \mreg/_08209_ ( .A(\mreg/_04251_ ), .ZN(\mreg/_02310_ ) );
OAI21_X1 \mreg/_08210_ ( .A(\mreg/_02309_ ), .B1(\mreg/_01374_ ), .B2(\mreg/_02310_ ), .ZN(\mreg/_02311_ ) );
AOI221_X4 \mreg/_08211_ ( .A(\mreg/_02311_ ), .B1(\mreg/_04187_ ), .B2(\mreg/_01465_ ), .C1(\mreg/_04155_ ), .C2(\mreg/_01505_ ), .ZN(\mreg/_02312_ ) );
AND4_X4 \mreg/_08212_ ( .A1(\mreg/_02300_ ), .A2(\mreg/_02304_ ), .A3(\mreg/_02308_ ), .A4(\mreg/_02312_ ), .ZN(\mreg/_02313_ ) );
AND3_X1 \mreg/_08213_ ( .A1(\mreg/_01107_ ), .A2(\mreg/_01118_ ), .A3(\mreg/_04283_ ), .ZN(\mreg/_02314_ ) );
AOI221_X4 \mreg/_08214_ ( .A(\mreg/_02314_ ), .B1(\mreg/_01219_ ), .B2(\mreg/_04731_ ), .C1(\mreg/_04635_ ), .C2(\mreg/_01222_ ), .ZN(\mreg/_02315_ ) );
NAND3_X1 \mreg/_08215_ ( .A1(\mreg/_01059_ ), .A2(\mreg/_01436_ ), .A3(\mreg/_04795_ ), .ZN(\mreg/_02316_ ) );
NAND3_X1 \mreg/_08216_ ( .A1(\mreg/_01092_ ), .A2(\mreg/_01282_ ), .A3(\mreg/_04827_ ), .ZN(\mreg/_02317_ ) );
NAND3_X1 \mreg/_08217_ ( .A1(\mreg/_01381_ ), .A2(\mreg/_01306_ ), .A3(\mreg/_04859_ ), .ZN(\mreg/_02318_ ) );
NAND3_X1 \mreg/_08218_ ( .A1(\mreg/_01339_ ), .A2(\mreg/_01087_ ), .A3(\mreg/_04763_ ), .ZN(\mreg/_02319_ ) );
AND4_X1 \mreg/_08219_ ( .A1(\mreg/_02316_ ), .A2(\mreg/_02317_ ), .A3(\mreg/_02318_ ), .A4(\mreg/_02319_ ), .ZN(\mreg/_02320_ ) );
NAND3_X1 \mreg/_08220_ ( .A1(\mreg/_01301_ ), .A2(\mreg/_01289_ ), .A3(\mreg/_04091_ ), .ZN(\mreg/_02321_ ) );
NAND3_X1 \mreg/_08221_ ( .A1(\mreg/_01121_ ), .A2(\mreg/_01130_ ), .A3(\mreg/_04923_ ), .ZN(\mreg/_02322_ ) );
NAND3_X1 \mreg/_08222_ ( .A1(\mreg/_01117_ ), .A2(\mreg/_01144_ ), .A3(\mreg/_03963_ ), .ZN(\mreg/_02323_ ) );
NAND3_X1 \mreg/_08223_ ( .A1(\mreg/_01126_ ), .A2(\mreg/_01162_ ), .A3(\mreg/_04891_ ), .ZN(\mreg/_02324_ ) );
NAND3_X1 \mreg/_08224_ ( .A1(\mreg/_01112_ ), .A2(\mreg/_01217_ ), .A3(\mreg/_03995_ ), .ZN(\mreg/_02325_ ) );
AND4_X1 \mreg/_08225_ ( .A1(\mreg/_02322_ ), .A2(\mreg/_02323_ ), .A3(\mreg/_02324_ ), .A4(\mreg/_02325_ ), .ZN(\mreg/_02326_ ) );
NAND3_X1 \mreg/_08226_ ( .A1(\mreg/_01308_ ), .A2(\mreg/_01295_ ), .A3(\mreg/_04123_ ), .ZN(\mreg/_02327_ ) );
AND3_X1 \mreg/_08227_ ( .A1(\mreg/_01148_ ), .A2(\mreg/_01622_ ), .A3(\mreg/_04059_ ), .ZN(\mreg/_02328_ ) );
AND3_X1 \mreg/_08228_ ( .A1(\mreg/_01338_ ), .A2(\mreg/_04027_ ), .A3(\mreg/_01151_ ), .ZN(\mreg/_02329_ ) );
NOR2_X1 \mreg/_08229_ ( .A1(\mreg/_02328_ ), .A2(\mreg/_02329_ ), .ZN(\mreg/_02330_ ) );
AND4_X1 \mreg/_08230_ ( .A1(\mreg/_02321_ ), .A2(\mreg/_02326_ ), .A3(\mreg/_02327_ ), .A4(\mreg/_02330_ ), .ZN(\mreg/_02331_ ) );
NAND4_X1 \mreg/_08231_ ( .A1(\mreg/_02313_ ), .A2(\mreg/_02315_ ), .A3(\mreg/_02320_ ), .A4(\mreg/_02331_ ), .ZN(\mreg/_03931_ ) );
AND3_X1 \mreg/_08232_ ( .A1(\mreg/_01058_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04349_ ), .ZN(\mreg/_02332_ ) );
AOI221_X4 \mreg/_08233_ ( .A(\mreg/_02332_ ), .B1(\mreg/_04317_ ), .B2(\mreg/_01377_ ), .C1(\mreg/_04669_ ), .C2(\mreg/_01175_ ), .ZN(\mreg/_02333_ ) );
AOI22_X1 \mreg/_08234_ ( .A1(\mreg/_04829_ ), .A2(\mreg/_01431_ ), .B1(\mreg/_01363_ ), .B2(\mreg/_04925_ ), .ZN(\mreg/_02334_ ) );
INV_X1 \mreg/_08235_ ( .A(\mreg/_00060_ ), .ZN(\mreg/_02335_ ) );
AOI22_X1 \mreg/_08236_ ( .A1(\mreg/_01361_ ), .A2(\mreg/_03965_ ), .B1(\mreg/_01173_ ), .B2(\mreg/_02335_ ), .ZN(\mreg/_02336_ ) );
AND3_X1 \mreg/_08237_ ( .A1(\mreg/_02333_ ), .A2(\mreg/_02334_ ), .A3(\mreg/_02336_ ), .ZN(\mreg/_02337_ ) );
NAND3_X1 \mreg/_08238_ ( .A1(\mreg/_01156_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04477_ ), .ZN(\mreg/_02338_ ) );
NAND3_X1 \mreg/_08239_ ( .A1(\mreg/_01082_ ), .A2(\mreg/_04573_ ), .A3(\mreg/_01151_ ), .ZN(\mreg/_02339_ ) );
NAND3_X1 \mreg/_08240_ ( .A1(\mreg/_01092_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04381_ ), .ZN(\mreg/_02340_ ) );
NAND3_X1 \mreg/_08241_ ( .A1(\mreg/_01064_ ), .A2(\mreg/_01114_ ), .A3(\mreg/_04637_ ), .ZN(\mreg/_02341_ ) );
NAND3_X1 \mreg/_08242_ ( .A1(\mreg/_01338_ ), .A2(\mreg/_04029_ ), .A3(\mreg/_01151_ ), .ZN(\mreg/_02342_ ) );
AND4_X1 \mreg/_08243_ ( .A1(\mreg/_02339_ ), .A2(\mreg/_02340_ ), .A3(\mreg/_02341_ ), .A4(\mreg/_02342_ ), .ZN(\mreg/_02343_ ) );
NAND3_X1 \mreg/_08244_ ( .A1(\mreg/_01383_ ), .A2(\mreg/_01302_ ), .A3(\mreg/_04285_ ), .ZN(\mreg/_02344_ ) );
AOI22_X1 \mreg/_08245_ ( .A1(\mreg/_01228_ ), .A2(\mreg/_04797_ ), .B1(\mreg/_01080_ ), .B2(\mreg/_04157_ ), .ZN(\mreg/_02345_ ) );
AND4_X1 \mreg/_08246_ ( .A1(\mreg/_02338_ ), .A2(\mreg/_02343_ ), .A3(\mreg/_02344_ ), .A4(\mreg/_02345_ ), .ZN(\mreg/_02346_ ) );
INV_X1 \mreg/_08247_ ( .A(\mreg/_04093_ ), .ZN(\mreg/_02347_ ) );
INV_X1 \mreg/_08248_ ( .A(\mreg/_03997_ ), .ZN(\mreg/_02348_ ) );
OAI22_X1 \mreg/_08249_ ( .A1(\mreg/_02347_ ), .A2(\mreg/_01393_ ), .B1(\mreg/_01396_ ), .B2(\mreg/_02348_ ), .ZN(\mreg/_02349_ ) );
NAND3_X1 \mreg/_08250_ ( .A1(\mreg/_01381_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04413_ ), .ZN(\mreg/_02350_ ) );
NAND3_X1 \mreg/_08251_ ( .A1(\mreg/_01304_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04605_ ), .ZN(\mreg/_02351_ ) );
NAND3_X1 \mreg/_08252_ ( .A1(\mreg/_01177_ ), .A2(\mreg/_04445_ ), .A3(\mreg/_01251_ ), .ZN(\mreg/_02352_ ) );
NAND3_X1 \mreg/_08253_ ( .A1(\mreg/_01621_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04189_ ), .ZN(\mreg/_02353_ ) );
NAND4_X1 \mreg/_08254_ ( .A1(\mreg/_02350_ ), .A2(\mreg/_02351_ ), .A3(\mreg/_02352_ ), .A4(\mreg/_02353_ ), .ZN(\mreg/_02354_ ) );
AND3_X1 \mreg/_08255_ ( .A1(\mreg/_01098_ ), .A2(\mreg/_01387_ ), .A3(\mreg/_04861_ ), .ZN(\mreg/_02355_ ) );
AND3_X1 \mreg/_08256_ ( .A1(\mreg/_01250_ ), .A2(\mreg/_04893_ ), .A3(\mreg/_01251_ ), .ZN(\mreg/_02356_ ) );
NOR4_X1 \mreg/_08257_ ( .A1(\mreg/_02349_ ), .A2(\mreg/_02354_ ), .A3(\mreg/_02355_ ), .A4(\mreg/_02356_ ), .ZN(\mreg/_02357_ ) );
NAND3_X1 \mreg/_08258_ ( .A1(\mreg/_01339_ ), .A2(\mreg/_01087_ ), .A3(\mreg/_04765_ ), .ZN(\mreg/_02358_ ) );
INV_X1 \mreg/_08259_ ( .A(\mreg/_04733_ ), .ZN(\mreg/_02359_ ) );
OAI21_X1 \mreg/_08260_ ( .A(\mreg/_02358_ ), .B1(\mreg/_01786_ ), .B2(\mreg/_02359_ ), .ZN(\mreg/_02360_ ) );
NAND4_X1 \mreg/_08261_ ( .A1(\mreg/_01667_ ), .A2(\mreg/_01251_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04509_ ), .ZN(\mreg/_02361_ ) );
INV_X1 \mreg/_08262_ ( .A(\mreg/_04541_ ), .ZN(\mreg/_02362_ ) );
OAI21_X1 \mreg/_08263_ ( .A(\mreg/_02361_ ), .B1(\mreg/_01191_ ), .B2(\mreg/_02362_ ), .ZN(\mreg/_02363_ ) );
NAND4_X1 \mreg/_08264_ ( .A1(\mreg/_01667_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04221_ ), .A4(\mreg/_01981_ ), .ZN(\mreg/_02364_ ) );
INV_X1 \mreg/_08265_ ( .A(\mreg/_04253_ ), .ZN(\mreg/_02365_ ) );
OAI21_X1 \mreg/_08266_ ( .A(\mreg/_02364_ ), .B1(\mreg/_01069_ ), .B2(\mreg/_02365_ ), .ZN(\mreg/_02366_ ) );
NAND3_X1 \mreg/_08267_ ( .A1(\mreg/_01238_ ), .A2(\mreg/_01248_ ), .A3(\mreg/_04125_ ), .ZN(\mreg/_02367_ ) );
INV_X1 \mreg/_08268_ ( .A(\mreg/_04061_ ), .ZN(\mreg/_02368_ ) );
OAI21_X1 \mreg/_08269_ ( .A(\mreg/_02367_ ), .B1(\mreg/_01791_ ), .B2(\mreg/_02368_ ), .ZN(\mreg/_02369_ ) );
NOR4_X1 \mreg/_08270_ ( .A1(\mreg/_02360_ ), .A2(\mreg/_02363_ ), .A3(\mreg/_02366_ ), .A4(\mreg/_02369_ ), .ZN(\mreg/_02370_ ) );
NAND4_X1 \mreg/_08271_ ( .A1(\mreg/_02337_ ), .A2(\mreg/_02346_ ), .A3(\mreg/_02357_ ), .A4(\mreg/_02370_ ), .ZN(\mreg/_03933_ ) );
NAND3_X1 \mreg/_08272_ ( .A1(\mreg/_01146_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04606_ ), .ZN(\mreg/_02371_ ) );
NAND3_X1 \mreg/_08273_ ( .A1(\mreg/_01255_ ), .A2(\mreg/_04574_ ), .A3(\mreg/_01150_ ), .ZN(\mreg/_02372_ ) );
NAND2_X1 \mreg/_08274_ ( .A1(\mreg/_02371_ ), .A2(\mreg/_02372_ ), .ZN(\mreg/_02373_ ) );
INV_X1 \mreg/_08275_ ( .A(\mreg/_00061_ ), .ZN(\mreg/_02374_ ) );
AOI221_X4 \mreg/_08276_ ( .A(\mreg/_02373_ ), .B1(\mreg/_02374_ ), .B2(\mreg/_01172_ ), .C1(\mreg/_04670_ ), .C2(\mreg/_01175_ ), .ZN(\mreg/_02375_ ) );
NAND4_X1 \mreg/_08277_ ( .A1(\mreg/_01269_ ), .A2(\mreg/_01366_ ), .A3(\mreg/_03877_ ), .A4(\mreg/_04510_ ), .ZN(\mreg/_02376_ ) );
INV_X1 \mreg/_08278_ ( .A(\mreg/_04542_ ), .ZN(\mreg/_02377_ ) );
OAI21_X1 \mreg/_08279_ ( .A(\mreg/_02376_ ), .B1(\mreg/_01190_ ), .B2(\mreg/_02377_ ), .ZN(\mreg/_02378_ ) );
AOI221_X4 \mreg/_08280_ ( .A(\mreg/_02378_ ), .B1(\mreg/_04478_ ), .B2(\mreg/_01195_ ), .C1(\mreg/_04446_ ), .C2(\mreg/_01660_ ), .ZN(\mreg/_02379_ ) );
NAND3_X1 \mreg/_08281_ ( .A1(\mreg/_01398_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04382_ ), .ZN(\mreg/_02380_ ) );
NAND3_X1 \mreg/_08282_ ( .A1(\mreg/_01096_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04414_ ), .ZN(\mreg/_02381_ ) );
NAND2_X1 \mreg/_08283_ ( .A1(\mreg/_02380_ ), .A2(\mreg/_02381_ ), .ZN(\mreg/_02382_ ) );
AOI221_X4 \mreg/_08284_ ( .A(\mreg/_02382_ ), .B1(\mreg/_04350_ ), .B2(\mreg/_01204_ ), .C1(\mreg/_04318_ ), .C2(\mreg/_01377_ ), .ZN(\mreg/_02383_ ) );
NAND4_X1 \mreg/_08285_ ( .A1(\mreg/_01365_ ), .A2(\mreg/_03877_ ), .A3(\mreg/_04222_ ), .A4(\mreg/_01372_ ), .ZN(\mreg/_02384_ ) );
INV_X1 \mreg/_08286_ ( .A(\mreg/_04254_ ), .ZN(\mreg/_02385_ ) );
OAI21_X1 \mreg/_08287_ ( .A(\mreg/_02384_ ), .B1(\mreg/_01374_ ), .B2(\mreg/_02385_ ), .ZN(\mreg/_02386_ ) );
AOI221_X4 \mreg/_08288_ ( .A(\mreg/_02386_ ), .B1(\mreg/_04190_ ), .B2(\mreg/_01074_ ), .C1(\mreg/_04158_ ), .C2(\mreg/_01505_ ), .ZN(\mreg/_02387_ ) );
AND4_X1 \mreg/_08289_ ( .A1(\mreg/_02375_ ), .A2(\mreg/_02379_ ), .A3(\mreg/_02383_ ), .A4(\mreg/_02387_ ), .ZN(\mreg/_02388_ ) );
NAND3_X1 \mreg/_08290_ ( .A1(\mreg/_01275_ ), .A2(\mreg/_01287_ ), .A3(\mreg/_04830_ ), .ZN(\mreg/_02389_ ) );
AOI22_X1 \mreg/_08291_ ( .A1(\mreg/_01284_ ), .A2(\mreg/_04798_ ), .B1(\mreg/_04766_ ), .B2(\mreg/_01230_ ), .ZN(\mreg/_02390_ ) );
NAND3_X1 \mreg/_08292_ ( .A1(\mreg/_01281_ ), .A2(\mreg/_01302_ ), .A3(\mreg/_04862_ ), .ZN(\mreg/_02391_ ) );
NAND3_X1 \mreg/_08293_ ( .A1(\mreg/_01621_ ), .A2(\mreg/_01622_ ), .A3(\mreg/_04286_ ), .ZN(\mreg/_02392_ ) );
NAND3_X1 \mreg/_08294_ ( .A1(\mreg/_01386_ ), .A2(\mreg/_01622_ ), .A3(\mreg/_04638_ ), .ZN(\mreg/_02393_ ) );
NAND3_X1 \mreg/_08295_ ( .A1(\mreg/_01067_ ), .A2(\mreg/_01130_ ), .A3(\mreg/_04734_ ), .ZN(\mreg/_02394_ ) );
AND3_X1 \mreg/_08296_ ( .A1(\mreg/_02392_ ), .A2(\mreg/_02393_ ), .A3(\mreg/_02394_ ), .ZN(\mreg/_02395_ ) );
AND4_X1 \mreg/_08297_ ( .A1(\mreg/_02389_ ), .A2(\mreg/_02390_ ), .A3(\mreg/_02391_ ), .A4(\mreg/_02395_ ), .ZN(\mreg/_02396_ ) );
NAND3_X1 \mreg/_08298_ ( .A1(\mreg/_01155_ ), .A2(\mreg/_01436_ ), .A3(\mreg/_04926_ ), .ZN(\mreg/_02397_ ) );
NAND3_X1 \mreg/_08299_ ( .A1(\mreg/_01158_ ), .A2(\mreg/_01282_ ), .A3(\mreg/_03966_ ), .ZN(\mreg/_02398_ ) );
NAND3_X1 \mreg/_08300_ ( .A1(\mreg/_01339_ ), .A2(\mreg/_01293_ ), .A3(\mreg/_04894_ ), .ZN(\mreg/_02399_ ) );
NAND3_X1 \mreg/_08301_ ( .A1(\mreg/_01113_ ), .A2(\mreg/_01477_ ), .A3(\mreg/_03998_ ), .ZN(\mreg/_02400_ ) );
AND4_X1 \mreg/_08302_ ( .A1(\mreg/_02397_ ), .A2(\mreg/_02398_ ), .A3(\mreg/_02399_ ), .A4(\mreg/_02400_ ), .ZN(\mreg/_02401_ ) );
AND3_X1 \mreg/_08303_ ( .A1(\mreg/_01232_ ), .A2(\mreg/_01233_ ), .A3(\mreg/_04094_ ), .ZN(\mreg/_02402_ ) );
AND3_X1 \mreg/_08304_ ( .A1(\mreg/_01304_ ), .A2(\mreg/_01384_ ), .A3(\mreg/_04062_ ), .ZN(\mreg/_02403_ ) );
AND3_X1 \mreg/_08305_ ( .A1(\mreg/_01238_ ), .A2(\mreg/_01248_ ), .A3(\mreg/_04126_ ), .ZN(\mreg/_02404_ ) );
AND3_X1 \mreg/_08306_ ( .A1(\mreg/_01291_ ), .A2(\mreg/_04030_ ), .A3(\mreg/_01391_ ), .ZN(\mreg/_02405_ ) );
NOR4_X1 \mreg/_08307_ ( .A1(\mreg/_02402_ ), .A2(\mreg/_02403_ ), .A3(\mreg/_02404_ ), .A4(\mreg/_02405_ ), .ZN(\mreg/_02406_ ) );
NAND4_X1 \mreg/_08308_ ( .A1(\mreg/_02388_ ), .A2(\mreg/_02396_ ), .A3(\mreg/_02401_ ), .A4(\mreg/_02406_ ), .ZN(\mreg/_03934_ ) );
NOR2_X4 \mreg/_08309_ ( .A1(\mreg/_03871_ ), .A2(\mreg/_03870_ ), .ZN(\mreg/_02407_ ) );
INV_X1 \mreg/_08310_ ( .A(\mreg/_03868_ ), .ZN(\mreg/_02408_ ) );
AND3_X2 \mreg/_08311_ ( .A1(\mreg/_02407_ ), .A2(\mreg/_03869_ ), .A3(\mreg/_02408_ ), .ZN(\mreg/_02409_ ) );
INV_X2 \mreg/_08312_ ( .A(\mreg/_03872_ ), .ZN(\mreg/_02410_ ) );
BUF_X2 \mreg/_08313_ ( .A(\mreg/_02410_ ), .Z(\mreg/_02411_ ) );
AND3_X1 \mreg/_08314_ ( .A1(\mreg/_02409_ ), .A2(\mreg/_04614_ ), .A3(\mreg/_02411_ ), .ZN(\mreg/_02412_ ) );
AND2_X4 \mreg/_08315_ ( .A1(\mreg/_03869_ ), .A2(\mreg/_03868_ ), .ZN(\mreg/_02413_ ) );
AND2_X4 \mreg/_08316_ ( .A1(\mreg/_02413_ ), .A2(\mreg/_02407_ ), .ZN(\mreg/_02414_ ) );
CLKBUF_X2 \mreg/_08317_ ( .A(\mreg/_02410_ ), .Z(\mreg/_02415_ ) );
AND2_X2 \mreg/_08318_ ( .A1(\mreg/_02414_ ), .A2(\mreg/_02415_ ), .ZN(\mreg/_02416_ ) );
INV_X32 \mreg/_08319_ ( .A(\mreg/_03869_ ), .ZN(\mreg/_02417_ ) );
AND3_X1 \mreg/_08320_ ( .A1(\mreg/_02407_ ), .A2(\mreg/_02417_ ), .A3(\mreg/_03868_ ), .ZN(\mreg/_02418_ ) );
BUF_X4 \mreg/_08321_ ( .A(\mreg/_02418_ ), .Z(\mreg/_02419_ ) );
AND2_X4 \mreg/_08322_ ( .A1(\mreg/_02419_ ), .A2(\mreg/_02410_ ), .ZN(\mreg/_02420_ ) );
BUF_X4 \mreg/_08323_ ( .A(\mreg/_02420_ ), .Z(\mreg/_02421_ ) );
AOI221_X4 \mreg/_08324_ ( .A(\mreg/_02412_ ), .B1(\mreg/_02416_ ), .B2(\mreg/_04710_ ), .C1(\mreg/_04262_ ), .C2(\mreg/_02421_ ), .ZN(\mreg/_02422_ ) );
AND2_X4 \mreg/_08325_ ( .A1(\mreg/_03871_ ), .A2(\mreg/_03870_ ), .ZN(\mreg/_02423_ ) );
AND2_X2 \mreg/_08326_ ( .A1(\mreg/_02413_ ), .A2(\mreg/_02423_ ), .ZN(\mreg/_02424_ ) );
BUF_X4 \mreg/_08327_ ( .A(\mreg/_02424_ ), .Z(\mreg/_02425_ ) );
BUF_X4 \mreg/_08328_ ( .A(\mreg/_02425_ ), .Z(\mreg/_02426_ ) );
BUF_X4 \mreg/_08329_ ( .A(\mreg/_02410_ ), .Z(\mreg/_02427_ ) );
BUF_X4 \mreg/_08330_ ( .A(\mreg/_02427_ ), .Z(\mreg/_02428_ ) );
NAND3_X1 \mreg/_08331_ ( .A1(\mreg/_02426_ ), .A2(\mreg/_04102_ ), .A3(\mreg/_02428_ ), .ZN(\mreg/_02429_ ) );
AND3_X1 \mreg/_08332_ ( .A1(\mreg/_02423_ ), .A2(\mreg/_03869_ ), .A3(\mreg/_02408_ ), .ZN(\mreg/_02430_ ) );
BUF_X4 \mreg/_08333_ ( .A(\mreg/_02430_ ), .Z(\mreg/_02431_ ) );
BUF_X4 \mreg/_08334_ ( .A(\mreg/_02431_ ), .Z(\mreg/_02432_ ) );
BUF_X4 \mreg/_08335_ ( .A(\mreg/_02410_ ), .Z(\mreg/_02433_ ) );
BUF_X4 \mreg/_08336_ ( .A(\mreg/_02433_ ), .Z(\mreg/_02434_ ) );
NAND3_X1 \mreg/_08337_ ( .A1(\mreg/_02432_ ), .A2(\mreg/_04070_ ), .A3(\mreg/_02434_ ), .ZN(\mreg/_02435_ ) );
NAND2_X4 \mreg/_08338_ ( .A1(\mreg/_02417_ ), .A2(\mreg/_03868_ ), .ZN(\mreg/_02436_ ) );
INV_X32 \mreg/_08339_ ( .A(\mreg/_03871_ ), .ZN(\mreg/_02437_ ) );
INV_X32 \mreg/_08340_ ( .A(\mreg/_03870_ ), .ZN(\mreg/_02438_ ) );
NOR3_X1 \mreg/_08341_ ( .A1(\mreg/_02436_ ), .A2(\mreg/_02437_ ), .A3(\mreg/_02438_ ), .ZN(\mreg/_02439_ ) );
BUF_X4 \mreg/_08342_ ( .A(\mreg/_02439_ ), .Z(\mreg/_02440_ ) );
BUF_X4 \mreg/_08343_ ( .A(\mreg/_02440_ ), .Z(\mreg/_02441_ ) );
NAND3_X1 \mreg/_08344_ ( .A1(\mreg/_02441_ ), .A2(\mreg/_04038_ ), .A3(\mreg/_02434_ ), .ZN(\mreg/_02442_ ) );
NOR3_X1 \mreg/_08345_ ( .A1(\mreg/_03872_ ), .A2(\mreg/_03869_ ), .A3(\mreg/_03868_ ), .ZN(\mreg/_02443_ ) );
BUF_X4 \mreg/_08346_ ( .A(\mreg/_02443_ ), .Z(\mreg/_02444_ ) );
BUF_X4 \mreg/_08347_ ( .A(\mreg/_02444_ ), .Z(\mreg/_02445_ ) );
BUF_X4 \mreg/_08348_ ( .A(\mreg/_02423_ ), .Z(\mreg/_02446_ ) );
BUF_X4 \mreg/_08349_ ( .A(\mreg/_02446_ ), .Z(\mreg/_02447_ ) );
BUF_X4 \mreg/_08350_ ( .A(\mreg/_02447_ ), .Z(\mreg/_02448_ ) );
NAND3_X1 \mreg/_08351_ ( .A1(\mreg/_02445_ ), .A2(\mreg/_04006_ ), .A3(\mreg/_02448_ ), .ZN(\mreg/_02449_ ) );
AND4_X1 \mreg/_08352_ ( .A1(\mreg/_02429_ ), .A2(\mreg/_02435_ ), .A3(\mreg/_02442_ ), .A4(\mreg/_02449_ ), .ZN(\mreg/_02450_ ) );
NOR2_X4 \mreg/_08353_ ( .A1(\mreg/_02417_ ), .A2(\mreg/_03868_ ), .ZN(\mreg/_02451_ ) );
NOR2_X1 \mreg/_08354_ ( .A1(\mreg/_02438_ ), .A2(\mreg/_03871_ ), .ZN(\mreg/_02452_ ) );
AND2_X2 \mreg/_08355_ ( .A1(\mreg/_02451_ ), .A2(\mreg/_02452_ ), .ZN(\mreg/_02453_ ) );
BUF_X4 \mreg/_08356_ ( .A(\mreg/_02453_ ), .Z(\mreg/_02454_ ) );
BUF_X4 \mreg/_08357_ ( .A(\mreg/_02454_ ), .Z(\mreg/_02455_ ) );
NAND3_X1 \mreg/_08358_ ( .A1(\mreg/_02455_ ), .A2(\mreg/_04806_ ), .A3(\mreg/_02428_ ), .ZN(\mreg/_02456_ ) );
AND3_X4 \mreg/_08359_ ( .A1(\mreg/_02413_ ), .A2(\mreg/_02437_ ), .A3(\mreg/_03870_ ), .ZN(\mreg/_02457_ ) );
BUF_X8 \mreg/_08360_ ( .A(\mreg/_02457_ ), .Z(\mreg/_02458_ ) );
BUF_X4 \mreg/_08361_ ( .A(\mreg/_02458_ ), .Z(\mreg/_02459_ ) );
BUF_X4 \mreg/_08362_ ( .A(\mreg/_02427_ ), .Z(\mreg/_02460_ ) );
NAND3_X1 \mreg/_08363_ ( .A1(\mreg/_02459_ ), .A2(\mreg/_04838_ ), .A3(\mreg/_02460_ ), .ZN(\mreg/_02461_ ) );
NOR3_X4 \mreg/_08364_ ( .A1(\mreg/_02436_ ), .A2(\mreg/_03871_ ), .A3(\mreg/_02438_ ), .ZN(\mreg/_02462_ ) );
BUF_X4 \mreg/_08365_ ( .A(\mreg/_02462_ ), .Z(\mreg/_02463_ ) );
BUF_X4 \mreg/_08366_ ( .A(\mreg/_02433_ ), .Z(\mreg/_02464_ ) );
NAND3_X1 \mreg/_08367_ ( .A1(\mreg/_02463_ ), .A2(\mreg/_04774_ ), .A3(\mreg/_02464_ ), .ZN(\mreg/_02465_ ) );
BUF_X4 \mreg/_08368_ ( .A(\mreg/_02452_ ), .Z(\mreg/_02466_ ) );
BUF_X2 \mreg/_08369_ ( .A(\mreg/_02466_ ), .Z(\mreg/_02467_ ) );
NAND3_X1 \mreg/_08370_ ( .A1(\mreg/_02445_ ), .A2(\mreg/_02467_ ), .A3(\mreg/_04742_ ), .ZN(\mreg/_02468_ ) );
AND4_X1 \mreg/_08371_ ( .A1(\mreg/_02456_ ), .A2(\mreg/_02461_ ), .A3(\mreg/_02465_ ), .A4(\mreg/_02468_ ), .ZN(\mreg/_02469_ ) );
NOR3_X1 \mreg/_08372_ ( .A1(\mreg/_02436_ ), .A2(\mreg/_02437_ ), .A3(\mreg/_03870_ ), .ZN(\mreg/_02470_ ) );
BUF_X4 \mreg/_08373_ ( .A(\mreg/_02470_ ), .Z(\mreg/_02471_ ) );
BUF_X4 \mreg/_08374_ ( .A(\mreg/_02471_ ), .Z(\mreg/_02472_ ) );
NAND3_X1 \mreg/_08375_ ( .A1(\mreg/_02472_ ), .A2(\mreg/_04902_ ), .A3(\mreg/_02428_ ), .ZN(\mreg/_02473_ ) );
NOR2_X4 \mreg/_08376_ ( .A1(\mreg/_02437_ ), .A2(\mreg/_03870_ ), .ZN(\mreg/_02474_ ) );
AND2_X1 \mreg/_08377_ ( .A1(\mreg/_02451_ ), .A2(\mreg/_02474_ ), .ZN(\mreg/_02475_ ) );
BUF_X4 \mreg/_08378_ ( .A(\mreg/_02475_ ), .Z(\mreg/_02476_ ) );
BUF_X4 \mreg/_08379_ ( .A(\mreg/_02476_ ), .Z(\mreg/_02477_ ) );
NAND3_X1 \mreg/_08380_ ( .A1(\mreg/_02477_ ), .A2(\mreg/_03942_ ), .A3(\mreg/_02464_ ), .ZN(\mreg/_02478_ ) );
BUF_X4 \mreg/_08381_ ( .A(\mreg/_02444_ ), .Z(\mreg/_02479_ ) );
BUF_X4 \mreg/_08382_ ( .A(\mreg/_02474_ ), .Z(\mreg/_02480_ ) );
BUF_X4 \mreg/_08383_ ( .A(\mreg/_02480_ ), .Z(\mreg/_02481_ ) );
NAND3_X1 \mreg/_08384_ ( .A1(\mreg/_02479_ ), .A2(\mreg/_02481_ ), .A3(\mreg/_04870_ ), .ZN(\mreg/_02482_ ) );
AND3_X4 \mreg/_08385_ ( .A1(\mreg/_02413_ ), .A2(\mreg/_03871_ ), .A3(\mreg/_02438_ ), .ZN(\mreg/_02483_ ) );
BUF_X8 \mreg/_08386_ ( .A(\mreg/_02483_ ), .Z(\mreg/_02484_ ) );
BUF_X4 \mreg/_08387_ ( .A(\mreg/_02484_ ), .Z(\mreg/_02485_ ) );
BUF_X4 \mreg/_08388_ ( .A(\mreg/_02433_ ), .Z(\mreg/_02486_ ) );
NAND3_X1 \mreg/_08389_ ( .A1(\mreg/_02485_ ), .A2(\mreg/_03974_ ), .A3(\mreg/_02486_ ), .ZN(\mreg/_02487_ ) );
AND4_X1 \mreg/_08390_ ( .A1(\mreg/_02473_ ), .A2(\mreg/_02478_ ), .A3(\mreg/_02482_ ), .A4(\mreg/_02487_ ), .ZN(\mreg/_02488_ ) );
AND4_X1 \mreg/_08391_ ( .A1(\mreg/_02422_ ), .A2(\mreg/_02450_ ), .A3(\mreg/_02469_ ), .A4(\mreg/_02488_ ), .ZN(\mreg/_02489_ ) );
BUF_X2 \mreg/_08392_ ( .A(\mreg/_02409_ ), .Z(\mreg/_02490_ ) );
NAND3_X1 \mreg/_08393_ ( .A1(\mreg/_02490_ ), .A2(\mreg/_04198_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02491_ ) );
NAND2_X4 \mreg/_08394_ ( .A1(\mreg/_02414_ ), .A2(\mreg/_03872_ ), .ZN(\mreg/_02492_ ) );
BUF_X4 \mreg/_08395_ ( .A(\mreg/_02492_ ), .Z(\mreg/_02493_ ) );
OAI21_X1 \mreg/_08396_ ( .A(\mreg/_02491_ ), .B1(\mreg/_02493_ ), .B2(\mreg/_01070_ ), .ZN(\mreg/_02494_ ) );
AND2_X2 \mreg/_08397_ ( .A1(\mreg/_02418_ ), .A2(\mreg/_03872_ ), .ZN(\mreg/_02495_ ) );
BUF_X4 \mreg/_08398_ ( .A(\mreg/_02495_ ), .Z(\mreg/_02496_ ) );
NOR2_X4 \mreg/_08399_ ( .A1(\mreg/_03869_ ), .A2(\mreg/_03868_ ), .ZN(\mreg/_02497_ ) );
AND2_X4 \mreg/_08400_ ( .A1(\mreg/_02497_ ), .A2(\mreg/_03872_ ), .ZN(\mreg/_02498_ ) );
BUF_X4 \mreg/_08401_ ( .A(\mreg/_02407_ ), .Z(\mreg/_02499_ ) );
AND2_X2 \mreg/_08402_ ( .A1(\mreg/_02498_ ), .A2(\mreg/_02499_ ), .ZN(\mreg/_02500_ ) );
BUF_X4 \mreg/_08403_ ( .A(\mreg/_02500_ ), .Z(\mreg/_02501_ ) );
AOI221_X4 \mreg/_08404_ ( .A(\mreg/_02494_ ), .B1(\mreg/_04166_ ), .B2(\mreg/_02496_ ), .C1(\mreg/_04134_ ), .C2(\mreg/_02501_ ), .ZN(\mreg/_02502_ ) );
BUF_X4 \mreg/_08405_ ( .A(\mreg/_02462_ ), .Z(\mreg/_02503_ ) );
BUF_X4 \mreg/_08406_ ( .A(\mreg/_02503_ ), .Z(\mreg/_02504_ ) );
NAND3_X1 \mreg/_08407_ ( .A1(\mreg/_02504_ ), .A2(\mreg/_04326_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02505_ ) );
BUF_X4 \mreg/_08408_ ( .A(\mreg/_02455_ ), .Z(\mreg/_02506_ ) );
NAND3_X1 \mreg/_08409_ ( .A1(\mreg/_02506_ ), .A2(\mreg/_04358_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02507_ ) );
BUF_X4 \mreg/_08410_ ( .A(\mreg/_02459_ ), .Z(\mreg/_02508_ ) );
NAND3_X1 \mreg/_08411_ ( .A1(\mreg/_02508_ ), .A2(\mreg/_04390_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02509_ ) );
BUF_X4 \mreg/_08412_ ( .A(\mreg/_02498_ ), .Z(\mreg/_02510_ ) );
BUF_X2 \mreg/_08413_ ( .A(\mreg/_02510_ ), .Z(\mreg/_02511_ ) );
BUF_X4 \mreg/_08414_ ( .A(\mreg/_02466_ ), .Z(\mreg/_02512_ ) );
BUF_X4 \mreg/_08415_ ( .A(\mreg/_02512_ ), .Z(\mreg/_02513_ ) );
NAND3_X1 \mreg/_08416_ ( .A1(\mreg/_02511_ ), .A2(\mreg/_04294_ ), .A3(\mreg/_02513_ ), .ZN(\mreg/_02514_ ) );
AND4_X1 \mreg/_08417_ ( .A1(\mreg/_02505_ ), .A2(\mreg/_02507_ ), .A3(\mreg/_02509_ ), .A4(\mreg/_02514_ ), .ZN(\mreg/_02515_ ) );
BUF_X4 \mreg/_08418_ ( .A(\mreg/_02432_ ), .Z(\mreg/_02516_ ) );
NAND3_X1 \mreg/_08419_ ( .A1(\mreg/_02516_ ), .A2(\mreg/_04646_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02517_ ) );
NAND3_X1 \mreg/_08420_ ( .A1(\mreg/_02472_ ), .A2(\mreg/_04454_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02518_ ) );
NAND3_X1 \mreg/_08421_ ( .A1(\mreg/_02477_ ), .A2(\mreg/_04486_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02519_ ) );
BUF_X2 \mreg/_08422_ ( .A(\mreg/_02510_ ), .Z(\mreg/_02520_ ) );
NAND3_X1 \mreg/_08423_ ( .A1(\mreg/_02520_ ), .A2(\mreg/_04422_ ), .A3(\mreg/_02481_ ), .ZN(\mreg/_02521_ ) );
NAND3_X1 \mreg/_08424_ ( .A1(\mreg/_02485_ ), .A2(\mreg/_04518_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02522_ ) );
AND4_X1 \mreg/_08425_ ( .A1(\mreg/_02518_ ), .A2(\mreg/_02519_ ), .A3(\mreg/_02521_ ), .A4(\mreg/_02522_ ), .ZN(\mreg/_02523_ ) );
BUF_X4 \mreg/_08426_ ( .A(\mreg/_02426_ ), .Z(\mreg/_02524_ ) );
NAND3_X1 \mreg/_08427_ ( .A1(\mreg/_02524_ ), .A2(\mreg/_04678_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02525_ ) );
AND3_X1 \mreg/_08428_ ( .A1(\mreg/_02520_ ), .A2(\mreg/_04550_ ), .A3(\mreg/_02447_ ), .ZN(\mreg/_02526_ ) );
AND2_X1 \mreg/_08429_ ( .A1(\mreg/_02440_ ), .A2(\mreg/_03872_ ), .ZN(\mreg/_02527_ ) );
AOI21_X1 \mreg/_08430_ ( .A(\mreg/_02526_ ), .B1(\mreg/_02527_ ), .B2(\mreg/_04582_ ), .ZN(\mreg/_02528_ ) );
AND4_X1 \mreg/_08431_ ( .A1(\mreg/_02517_ ), .A2(\mreg/_02523_ ), .A3(\mreg/_02525_ ), .A4(\mreg/_02528_ ), .ZN(\mreg/_02529_ ) );
NAND4_X1 \mreg/_08432_ ( .A1(\mreg/_02489_ ), .A2(\mreg/_02502_ ), .A3(\mreg/_02515_ ), .A4(\mreg/_02529_ ), .ZN(\mreg/_03878_ ) );
BUF_X4 \mreg/_08433_ ( .A(\mreg/_02510_ ), .Z(\mreg/_02530_ ) );
BUF_X4 \mreg/_08434_ ( .A(\mreg/_02530_ ), .Z(\mreg/_02531_ ) );
BUF_X4 \mreg/_08435_ ( .A(\mreg/_02447_ ), .Z(\mreg/_02532_ ) );
BUF_X4 \mreg/_08436_ ( .A(\mreg/_02532_ ), .Z(\mreg/_02533_ ) );
NAND3_X1 \mreg/_08437_ ( .A1(\mreg/_02531_ ), .A2(\mreg/_04561_ ), .A3(\mreg/_02533_ ), .ZN(\mreg/_02534_ ) );
BUF_X4 \mreg/_08438_ ( .A(\mreg/_02451_ ), .Z(\mreg/_02535_ ) );
BUF_X2 \mreg/_08439_ ( .A(\mreg/_02474_ ), .Z(\mreg/_02536_ ) );
NAND4_X1 \mreg/_08440_ ( .A1(\mreg/_02535_ ), .A2(\mreg/_02536_ ), .A3(\mreg/_04497_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_02537_ ) );
NAND2_X4 \mreg/_08441_ ( .A1(\mreg/_02484_ ), .A2(\mreg/_03872_ ), .ZN(\mreg/_02538_ ) );
BUF_X8 \mreg/_08442_ ( .A(\mreg/_02538_ ), .Z(\mreg/_02539_ ) );
OAI21_X1 \mreg/_08443_ ( .A(\mreg/_02537_ ), .B1(\mreg/_02539_ ), .B2(\mreg/_01192_ ), .ZN(\mreg/_02540_ ) );
AND2_X2 \mreg/_08444_ ( .A1(\mreg/_02470_ ), .A2(\mreg/_03872_ ), .ZN(\mreg/_02541_ ) );
BUF_X4 \mreg/_08445_ ( .A(\mreg/_02541_ ), .Z(\mreg/_02542_ ) );
AND2_X2 \mreg/_08446_ ( .A1(\mreg/_02498_ ), .A2(\mreg/_02474_ ), .ZN(\mreg/_02543_ ) );
BUF_X4 \mreg/_08447_ ( .A(\mreg/_02543_ ), .Z(\mreg/_02544_ ) );
AOI221_X4 \mreg/_08448_ ( .A(\mreg/_02540_ ), .B1(\mreg/_04465_ ), .B2(\mreg/_02542_ ), .C1(\mreg/_04433_ ), .C2(\mreg/_02544_ ), .ZN(\mreg/_02545_ ) );
BUF_X4 \mreg/_08449_ ( .A(\mreg/_02441_ ), .Z(\mreg/_02546_ ) );
NAND3_X1 \mreg/_08450_ ( .A1(\mreg/_02546_ ), .A2(\mreg/_04593_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02547_ ) );
AND3_X1 \mreg/_08451_ ( .A1(\mreg/_02432_ ), .A2(\mreg/_04657_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02548_ ) );
AND2_X2 \mreg/_08452_ ( .A1(\mreg/_02424_ ), .A2(\mreg/_03872_ ), .ZN(\mreg/_02549_ ) );
BUF_X4 \mreg/_08453_ ( .A(\mreg/_02549_ ), .Z(\mreg/_02550_ ) );
AOI21_X1 \mreg/_08454_ ( .A(\mreg/_02548_ ), .B1(\mreg/_01185_ ), .B2(\mreg/_02550_ ), .ZN(\mreg/_02551_ ) );
AND4_X4 \mreg/_08455_ ( .A1(\mreg/_02534_ ), .A2(\mreg/_02545_ ), .A3(\mreg/_02547_ ), .A4(\mreg/_02551_ ), .ZN(\mreg/_02552_ ) );
BUF_X2 \mreg/_08456_ ( .A(\mreg/_02410_ ), .Z(\mreg/_02553_ ) );
AND3_X1 \mreg/_08457_ ( .A1(\mreg/_02409_ ), .A2(\mreg/_04625_ ), .A3(\mreg/_02553_ ), .ZN(\mreg/_02554_ ) );
AOI221_X4 \mreg/_08458_ ( .A(\mreg/_02554_ ), .B1(\mreg/_02416_ ), .B2(\mreg/_04721_ ), .C1(\mreg/_04273_ ), .C2(\mreg/_02421_ ), .ZN(\mreg/_02555_ ) );
AND3_X1 \mreg/_08459_ ( .A1(\mreg/_02484_ ), .A2(\mreg/_03985_ ), .A3(\mreg/_02553_ ), .ZN(\mreg/_02556_ ) );
NAND3_X1 \mreg/_08460_ ( .A1(\mreg/_02471_ ), .A2(\mreg/_04913_ ), .A3(\mreg/_02411_ ), .ZN(\mreg/_02557_ ) );
NAND3_X1 \mreg/_08461_ ( .A1(\mreg/_02443_ ), .A2(\mreg/_02480_ ), .A3(\mreg/_04881_ ), .ZN(\mreg/_02558_ ) );
NAND2_X1 \mreg/_08462_ ( .A1(\mreg/_02557_ ), .A2(\mreg/_02558_ ), .ZN(\mreg/_02559_ ) );
AND2_X2 \mreg/_08463_ ( .A1(\mreg/_02476_ ), .A2(\mreg/_02415_ ), .ZN(\mreg/_02560_ ) );
AOI211_X4 \mreg/_08464_ ( .A(\mreg/_02556_ ), .B(\mreg/_02559_ ), .C1(\mreg/_03953_ ), .C2(\mreg/_02560_ ), .ZN(\mreg/_02561_ ) );
NAND3_X1 \mreg/_08465_ ( .A1(\mreg/_02463_ ), .A2(\mreg/_04785_ ), .A3(\mreg/_02434_ ), .ZN(\mreg/_02562_ ) );
BUF_X2 \mreg/_08466_ ( .A(\mreg/_02433_ ), .Z(\mreg/_02563_ ) );
NAND3_X1 \mreg/_08467_ ( .A1(\mreg/_02454_ ), .A2(\mreg/_04817_ ), .A3(\mreg/_02563_ ), .ZN(\mreg/_02564_ ) );
BUF_X2 \mreg/_08468_ ( .A(\mreg/_02458_ ), .Z(\mreg/_02565_ ) );
BUF_X2 \mreg/_08469_ ( .A(\mreg/_02433_ ), .Z(\mreg/_02566_ ) );
NAND3_X1 \mreg/_08470_ ( .A1(\mreg/_02565_ ), .A2(\mreg/_04849_ ), .A3(\mreg/_02566_ ), .ZN(\mreg/_02567_ ) );
BUF_X2 \mreg/_08471_ ( .A(\mreg/_02452_ ), .Z(\mreg/_02568_ ) );
NAND3_X1 \mreg/_08472_ ( .A1(\mreg/_02479_ ), .A2(\mreg/_02568_ ), .A3(\mreg/_04753_ ), .ZN(\mreg/_02569_ ) );
AND4_X1 \mreg/_08473_ ( .A1(\mreg/_02562_ ), .A2(\mreg/_02564_ ), .A3(\mreg/_02567_ ), .A4(\mreg/_02569_ ), .ZN(\mreg/_02570_ ) );
BUF_X2 \mreg/_08474_ ( .A(\mreg/_02431_ ), .Z(\mreg/_02571_ ) );
BUF_X2 \mreg/_08475_ ( .A(\mreg/_02411_ ), .Z(\mreg/_02572_ ) );
AND3_X1 \mreg/_08476_ ( .A1(\mreg/_02571_ ), .A2(\mreg/_04081_ ), .A3(\mreg/_02572_ ), .ZN(\mreg/_02573_ ) );
AND3_X1 \mreg/_08477_ ( .A1(\mreg/_02440_ ), .A2(\mreg/_04049_ ), .A3(\mreg/_02427_ ), .ZN(\mreg/_02574_ ) );
AND3_X1 \mreg/_08478_ ( .A1(\mreg/_02425_ ), .A2(\mreg/_04113_ ), .A3(\mreg/_02427_ ), .ZN(\mreg/_02575_ ) );
AND3_X1 \mreg/_08479_ ( .A1(\mreg/_02444_ ), .A2(\mreg/_04017_ ), .A3(\mreg/_02447_ ), .ZN(\mreg/_02576_ ) );
NOR4_X1 \mreg/_08480_ ( .A1(\mreg/_02573_ ), .A2(\mreg/_02574_ ), .A3(\mreg/_02575_ ), .A4(\mreg/_02576_ ), .ZN(\mreg/_02577_ ) );
AND4_X1 \mreg/_08481_ ( .A1(\mreg/_02555_ ), .A2(\mreg/_02561_ ), .A3(\mreg/_02570_ ), .A4(\mreg/_02577_ ), .ZN(\mreg/_02578_ ) );
BUF_X4 \mreg/_08482_ ( .A(\mreg/_02499_ ), .Z(\mreg/_02579_ ) );
BUF_X4 \mreg/_08483_ ( .A(\mreg/_02579_ ), .Z(\mreg/_02580_ ) );
BUF_X4 \mreg/_08484_ ( .A(\mreg/_02580_ ), .Z(\mreg/_02581_ ) );
NAND3_X1 \mreg/_08485_ ( .A1(\mreg/_02531_ ), .A2(\mreg/_04145_ ), .A3(\mreg/_02581_ ), .ZN(\mreg/_02582_ ) );
BUF_X4 \mreg/_08486_ ( .A(\mreg/_02419_ ), .Z(\mreg/_02583_ ) );
NAND3_X1 \mreg/_08487_ ( .A1(\mreg/_02583_ ), .A2(\mreg/_04177_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02584_ ) );
BUF_X4 \mreg/_08488_ ( .A(\mreg/_02451_ ), .Z(\mreg/_02585_ ) );
BUF_X4 \mreg/_08489_ ( .A(\mreg/_02585_ ), .Z(\mreg/_02586_ ) );
BUF_X4 \mreg/_08490_ ( .A(\mreg/_02586_ ), .Z(\mreg/_02587_ ) );
NAND4_X1 \mreg/_08491_ ( .A1(\mreg/_02587_ ), .A2(\mreg/_04209_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02581_ ), .ZN(\mreg/_02588_ ) );
BUF_X2 \mreg/_08492_ ( .A(\mreg/_02413_ ), .Z(\mreg/_02589_ ) );
NAND4_X1 \mreg/_08493_ ( .A1(\mreg/_02589_ ), .A2(\mreg/_02581_ ), .A3(\mreg/_04241_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_02590_ ) );
AND4_X1 \mreg/_08494_ ( .A1(\mreg/_02582_ ), .A2(\mreg/_02584_ ), .A3(\mreg/_02588_ ), .A4(\mreg/_02590_ ), .ZN(\mreg/_02591_ ) );
NAND3_X1 \mreg/_08495_ ( .A1(\mreg/_02506_ ), .A2(\mreg/_04369_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02592_ ) );
NAND3_X1 \mreg/_08496_ ( .A1(\mreg/_02508_ ), .A2(\mreg/_04401_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02593_ ) );
NAND3_X1 \mreg/_08497_ ( .A1(\mreg/_02503_ ), .A2(\mreg/_04337_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02594_ ) );
NAND3_X1 \mreg/_08498_ ( .A1(\mreg/_02511_ ), .A2(\mreg/_04305_ ), .A3(\mreg/_02513_ ), .ZN(\mreg/_02595_ ) );
AND4_X1 \mreg/_08499_ ( .A1(\mreg/_02592_ ), .A2(\mreg/_02593_ ), .A3(\mreg/_02594_ ), .A4(\mreg/_02595_ ), .ZN(\mreg/_02596_ ) );
NAND4_X1 \mreg/_08500_ ( .A1(\mreg/_02552_ ), .A2(\mreg/_02578_ ), .A3(\mreg/_02591_ ), .A4(\mreg/_02596_ ), .ZN(\mreg/_03889_ ) );
BUF_X4 \mreg/_08501_ ( .A(\mreg/_02439_ ), .Z(\mreg/_02597_ ) );
NAND3_X1 \mreg/_08502_ ( .A1(\mreg/_02597_ ), .A2(\mreg/_04604_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02598_ ) );
BUF_X2 \mreg/_08503_ ( .A(\mreg/_02498_ ), .Z(\mreg/_02599_ ) );
NAND3_X1 \mreg/_08504_ ( .A1(\mreg/_02599_ ), .A2(\mreg/_04572_ ), .A3(\mreg/_02446_ ), .ZN(\mreg/_02600_ ) );
NAND2_X1 \mreg/_08505_ ( .A1(\mreg/_02598_ ), .A2(\mreg/_02600_ ), .ZN(\mreg/_02601_ ) );
AND2_X1 \mreg/_08506_ ( .A1(\mreg/_02430_ ), .A2(\mreg/_03872_ ), .ZN(\mreg/_02602_ ) );
BUF_X4 \mreg/_08507_ ( .A(\mreg/_02602_ ), .Z(\mreg/_02603_ ) );
AOI221_X4 \mreg/_08508_ ( .A(\mreg/_02601_ ), .B1(\mreg/_01258_ ), .B2(\mreg/_02550_ ), .C1(\mreg/_04668_ ), .C2(\mreg/_02603_ ), .ZN(\mreg/_02604_ ) );
NAND4_X1 \mreg/_08509_ ( .A1(\mreg/_02535_ ), .A2(\mreg/_02536_ ), .A3(\mreg/_04508_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_02605_ ) );
OAI21_X1 \mreg/_08510_ ( .A(\mreg/_02605_ ), .B1(\mreg/_02539_ ), .B2(\mreg/_01262_ ), .ZN(\mreg/_02606_ ) );
AOI221_X4 \mreg/_08511_ ( .A(\mreg/_02606_ ), .B1(\mreg/_04476_ ), .B2(\mreg/_02542_ ), .C1(\mreg/_04444_ ), .C2(\mreg/_02544_ ), .ZN(\mreg/_02607_ ) );
BUF_X4 \mreg/_08512_ ( .A(\mreg/_02451_ ), .Z(\mreg/_02608_ ) );
BUF_X4 \mreg/_08513_ ( .A(\mreg/_02407_ ), .Z(\mreg/_02609_ ) );
NAND4_X1 \mreg/_08514_ ( .A1(\mreg/_02608_ ), .A2(\mreg/_04220_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02609_ ), .ZN(\mreg/_02610_ ) );
BUF_X4 \mreg/_08515_ ( .A(\mreg/_02492_ ), .Z(\mreg/_02611_ ) );
OAI21_X1 \mreg/_08516_ ( .A(\mreg/_02610_ ), .B1(\mreg/_02611_ ), .B2(\mreg/_01271_ ), .ZN(\mreg/_02612_ ) );
BUF_X4 \mreg/_08517_ ( .A(\mreg/_02495_ ), .Z(\mreg/_02613_ ) );
BUF_X4 \mreg/_08518_ ( .A(\mreg/_02500_ ), .Z(\mreg/_02614_ ) );
AOI221_X4 \mreg/_08519_ ( .A(\mreg/_02612_ ), .B1(\mreg/_04188_ ), .B2(\mreg/_02613_ ), .C1(\mreg/_04156_ ), .C2(\mreg/_02614_ ), .ZN(\mreg/_02615_ ) );
NAND3_X1 \mreg/_08520_ ( .A1(\mreg/_02455_ ), .A2(\mreg/_04380_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02616_ ) );
NAND3_X1 \mreg/_08521_ ( .A1(\mreg/_02459_ ), .A2(\mreg/_04412_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02617_ ) );
NAND3_X1 \mreg/_08522_ ( .A1(\mreg/_02463_ ), .A2(\mreg/_04348_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02618_ ) );
CLKBUF_X2 \mreg/_08523_ ( .A(\mreg/_02510_ ), .Z(\mreg/_02619_ ) );
NAND3_X1 \mreg/_08524_ ( .A1(\mreg/_02619_ ), .A2(\mreg/_04316_ ), .A3(\mreg/_02467_ ), .ZN(\mreg/_02620_ ) );
AND4_X1 \mreg/_08525_ ( .A1(\mreg/_02616_ ), .A2(\mreg/_02617_ ), .A3(\mreg/_02618_ ), .A4(\mreg/_02620_ ), .ZN(\mreg/_02621_ ) );
AND4_X2 \mreg/_08526_ ( .A1(\mreg/_02604_ ), .A2(\mreg/_02607_ ), .A3(\mreg/_02615_ ), .A4(\mreg/_02621_ ), .ZN(\mreg/_02622_ ) );
BUF_X4 \mreg/_08527_ ( .A(\mreg/_02427_ ), .Z(\mreg/_02623_ ) );
BUF_X4 \mreg/_08528_ ( .A(\mreg/_02623_ ), .Z(\mreg/_02624_ ) );
NAND3_X1 \mreg/_08529_ ( .A1(\mreg/_02504_ ), .A2(\mreg/_04796_ ), .A3(\mreg/_02624_ ), .ZN(\mreg/_02625_ ) );
AND3_X1 \mreg/_08530_ ( .A1(\mreg/_02414_ ), .A2(\mreg/_04732_ ), .A3(\mreg/_02415_ ), .ZN(\mreg/_02626_ ) );
AND2_X2 \mreg/_08531_ ( .A1(\mreg/_02409_ ), .A2(\mreg/_02410_ ), .ZN(\mreg/_02627_ ) );
AOI221_X4 \mreg/_08532_ ( .A(\mreg/_02626_ ), .B1(\mreg/_02627_ ), .B2(\mreg/_04636_ ), .C1(\mreg/_04284_ ), .C2(\mreg/_02420_ ), .ZN(\mreg/_02628_ ) );
BUF_X4 \mreg/_08533_ ( .A(\mreg/_02444_ ), .Z(\mreg/_02629_ ) );
BUF_X4 \mreg/_08534_ ( .A(\mreg/_02629_ ), .Z(\mreg/_02630_ ) );
NAND3_X1 \mreg/_08535_ ( .A1(\mreg/_02630_ ), .A2(\mreg/_02513_ ), .A3(\mreg/_04764_ ), .ZN(\mreg/_02631_ ) );
BUF_X2 \mreg/_08536_ ( .A(\mreg/_02458_ ), .Z(\mreg/_02632_ ) );
BUF_X2 \mreg/_08537_ ( .A(\mreg/_02411_ ), .Z(\mreg/_02633_ ) );
AND3_X1 \mreg/_08538_ ( .A1(\mreg/_02632_ ), .A2(\mreg/_04860_ ), .A3(\mreg/_02633_ ), .ZN(\mreg/_02634_ ) );
AND2_X2 \mreg/_08539_ ( .A1(\mreg/_02453_ ), .A2(\mreg/_02411_ ), .ZN(\mreg/_02635_ ) );
BUF_X4 \mreg/_08540_ ( .A(\mreg/_02635_ ), .Z(\mreg/_02636_ ) );
AOI21_X1 \mreg/_08541_ ( .A(\mreg/_02634_ ), .B1(\mreg/_04828_ ), .B2(\mreg/_02636_ ), .ZN(\mreg/_02637_ ) );
AND4_X1 \mreg/_08542_ ( .A1(\mreg/_02625_ ), .A2(\mreg/_02628_ ), .A3(\mreg/_02631_ ), .A4(\mreg/_02637_ ), .ZN(\mreg/_02638_ ) );
BUF_X2 \mreg/_08543_ ( .A(\mreg/_02471_ ), .Z(\mreg/_02639_ ) );
NAND3_X1 \mreg/_08544_ ( .A1(\mreg/_02639_ ), .A2(\mreg/_04924_ ), .A3(\mreg/_02624_ ), .ZN(\mreg/_02640_ ) );
BUF_X4 \mreg/_08545_ ( .A(\mreg/_02477_ ), .Z(\mreg/_02641_ ) );
BUF_X4 \mreg/_08546_ ( .A(\mreg/_02623_ ), .Z(\mreg/_02642_ ) );
NAND3_X1 \mreg/_08547_ ( .A1(\mreg/_02641_ ), .A2(\mreg/_03964_ ), .A3(\mreg/_02642_ ), .ZN(\mreg/_02643_ ) );
BUF_X2 \mreg/_08548_ ( .A(\mreg/_02536_ ), .Z(\mreg/_02644_ ) );
BUF_X2 \mreg/_08549_ ( .A(\mreg/_02644_ ), .Z(\mreg/_02645_ ) );
NAND3_X1 \mreg/_08550_ ( .A1(\mreg/_02630_ ), .A2(\mreg/_02645_ ), .A3(\mreg/_04892_ ), .ZN(\mreg/_02646_ ) );
BUF_X4 \mreg/_08551_ ( .A(\mreg/_02485_ ), .Z(\mreg/_02647_ ) );
BUF_X4 \mreg/_08552_ ( .A(\mreg/_02428_ ), .Z(\mreg/_02648_ ) );
NAND3_X1 \mreg/_08553_ ( .A1(\mreg/_02647_ ), .A2(\mreg/_03996_ ), .A3(\mreg/_02648_ ), .ZN(\mreg/_02649_ ) );
AND4_X1 \mreg/_08554_ ( .A1(\mreg/_02640_ ), .A2(\mreg/_02643_ ), .A3(\mreg/_02646_ ), .A4(\mreg/_02649_ ), .ZN(\mreg/_02650_ ) );
NAND3_X1 \mreg/_08555_ ( .A1(\mreg/_02630_ ), .A2(\mreg/_04028_ ), .A3(\mreg/_02533_ ), .ZN(\mreg/_02651_ ) );
BUF_X4 \mreg/_08556_ ( .A(\mreg/_02623_ ), .Z(\mreg/_02652_ ) );
NAND3_X1 \mreg/_08557_ ( .A1(\mreg/_02516_ ), .A2(\mreg/_04092_ ), .A3(\mreg/_02652_ ), .ZN(\mreg/_02653_ ) );
BUF_X4 \mreg/_08558_ ( .A(\mreg/_02623_ ), .Z(\mreg/_02654_ ) );
NAND3_X1 \mreg/_08559_ ( .A1(\mreg/_02546_ ), .A2(\mreg/_04060_ ), .A3(\mreg/_02654_ ), .ZN(\mreg/_02655_ ) );
NAND3_X1 \mreg/_08560_ ( .A1(\mreg/_02524_ ), .A2(\mreg/_04124_ ), .A3(\mreg/_02648_ ), .ZN(\mreg/_02656_ ) );
AND4_X1 \mreg/_08561_ ( .A1(\mreg/_02651_ ), .A2(\mreg/_02653_ ), .A3(\mreg/_02655_ ), .A4(\mreg/_02656_ ), .ZN(\mreg/_02657_ ) );
NAND4_X1 \mreg/_08562_ ( .A1(\mreg/_02622_ ), .A2(\mreg/_02638_ ), .A3(\mreg/_02650_ ), .A4(\mreg/_02657_ ), .ZN(\mreg/_03900_ ) );
NAND3_X1 \mreg/_08563_ ( .A1(\mreg/_02516_ ), .A2(\mreg/_04671_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02658_ ) );
NAND4_X1 \mreg/_08564_ ( .A1(\mreg/_02535_ ), .A2(\mreg/_02536_ ), .A3(\mreg/_04511_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_02659_ ) );
BUF_X4 \mreg/_08565_ ( .A(\mreg/_02538_ ), .Z(\mreg/_02660_ ) );
OAI21_X1 \mreg/_08566_ ( .A(\mreg/_02659_ ), .B1(\mreg/_02660_ ), .B2(\mreg/_01320_ ), .ZN(\mreg/_02661_ ) );
AOI221_X4 \mreg/_08567_ ( .A(\mreg/_02661_ ), .B1(\mreg/_04479_ ), .B2(\mreg/_02542_ ), .C1(\mreg/_04447_ ), .C2(\mreg/_02544_ ), .ZN(\mreg/_02662_ ) );
NAND3_X1 \mreg/_08568_ ( .A1(\mreg/_02524_ ), .A2(\mreg/_01315_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02663_ ) );
BUF_X2 \mreg/_08569_ ( .A(\mreg/_02447_ ), .Z(\mreg/_02664_ ) );
AND3_X1 \mreg/_08570_ ( .A1(\mreg/_02619_ ), .A2(\mreg/_04575_ ), .A3(\mreg/_02664_ ), .ZN(\mreg/_02665_ ) );
AOI21_X1 \mreg/_08571_ ( .A(\mreg/_02665_ ), .B1(\mreg/_02527_ ), .B2(\mreg/_04607_ ), .ZN(\mreg/_02666_ ) );
AND4_X4 \mreg/_08572_ ( .A1(\mreg/_02658_ ), .A2(\mreg/_02662_ ), .A3(\mreg/_02663_ ), .A4(\mreg/_02666_ ), .ZN(\mreg/_02667_ ) );
NAND4_X1 \mreg/_08573_ ( .A1(\mreg/_02586_ ), .A2(\mreg/_04223_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02580_ ), .ZN(\mreg/_02668_ ) );
NAND4_X1 \mreg/_08574_ ( .A1(\mreg/_02589_ ), .A2(\mreg/_02580_ ), .A3(\mreg/_04255_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_02669_ ) );
NAND2_X1 \mreg/_08575_ ( .A1(\mreg/_02668_ ), .A2(\mreg/_02669_ ), .ZN(\mreg/_02670_ ) );
AOI221_X4 \mreg/_08576_ ( .A(\mreg/_02670_ ), .B1(\mreg/_04191_ ), .B2(\mreg/_02496_ ), .C1(\mreg/_04159_ ), .C2(\mreg/_02501_ ), .ZN(\mreg/_02671_ ) );
BUF_X4 \mreg/_08577_ ( .A(\mreg/_02455_ ), .Z(\mreg/_02672_ ) );
NAND3_X1 \mreg/_08578_ ( .A1(\mreg/_02672_ ), .A2(\mreg/_04383_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02673_ ) );
BUF_X4 \mreg/_08579_ ( .A(\mreg/_02459_ ), .Z(\mreg/_02674_ ) );
NAND3_X1 \mreg/_08580_ ( .A1(\mreg/_02674_ ), .A2(\mreg/_04415_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02675_ ) );
NAND3_X1 \mreg/_08581_ ( .A1(\mreg/_02504_ ), .A2(\mreg/_04351_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02676_ ) );
NAND3_X1 \mreg/_08582_ ( .A1(\mreg/_02511_ ), .A2(\mreg/_04319_ ), .A3(\mreg/_02513_ ), .ZN(\mreg/_02677_ ) );
AND4_X1 \mreg/_08583_ ( .A1(\mreg/_02673_ ), .A2(\mreg/_02675_ ), .A3(\mreg/_02676_ ), .A4(\mreg/_02677_ ), .ZN(\mreg/_02678_ ) );
AND3_X1 \mreg/_08584_ ( .A1(\mreg/_02409_ ), .A2(\mreg/_04639_ ), .A3(\mreg/_02415_ ), .ZN(\mreg/_02679_ ) );
AOI221_X4 \mreg/_08585_ ( .A(\mreg/_02679_ ), .B1(\mreg/_02416_ ), .B2(\mreg/_04735_ ), .C1(\mreg/_04287_ ), .C2(\mreg/_02421_ ), .ZN(\mreg/_02680_ ) );
NAND3_X1 \mreg/_08586_ ( .A1(\mreg/_02463_ ), .A2(\mreg/_04799_ ), .A3(\mreg/_02460_ ), .ZN(\mreg/_02681_ ) );
NAND3_X1 \mreg/_08587_ ( .A1(\mreg/_02454_ ), .A2(\mreg/_04831_ ), .A3(\mreg/_02486_ ), .ZN(\mreg/_02682_ ) );
NAND3_X1 \mreg/_08588_ ( .A1(\mreg/_02632_ ), .A2(\mreg/_04863_ ), .A3(\mreg/_02572_ ), .ZN(\mreg/_02683_ ) );
BUF_X4 \mreg/_08589_ ( .A(\mreg/_02444_ ), .Z(\mreg/_02684_ ) );
NAND3_X1 \mreg/_08590_ ( .A1(\mreg/_02684_ ), .A2(\mreg/_02568_ ), .A3(\mreg/_04767_ ), .ZN(\mreg/_02685_ ) );
AND4_X1 \mreg/_08591_ ( .A1(\mreg/_02681_ ), .A2(\mreg/_02682_ ), .A3(\mreg/_02683_ ), .A4(\mreg/_02685_ ), .ZN(\mreg/_02686_ ) );
NAND3_X1 \mreg/_08592_ ( .A1(\mreg/_02471_ ), .A2(\mreg/_04927_ ), .A3(\mreg/_02464_ ), .ZN(\mreg/_02687_ ) );
BUF_X4 \mreg/_08593_ ( .A(\mreg/_02433_ ), .Z(\mreg/_02688_ ) );
NAND3_X1 \mreg/_08594_ ( .A1(\mreg/_02476_ ), .A2(\mreg/_03967_ ), .A3(\mreg/_02688_ ), .ZN(\mreg/_02689_ ) );
NAND3_X1 \mreg/_08595_ ( .A1(\mreg/_02684_ ), .A2(\mreg/_02481_ ), .A3(\mreg/_04895_ ), .ZN(\mreg/_02690_ ) );
BUF_X4 \mreg/_08596_ ( .A(\mreg/_02433_ ), .Z(\mreg/_02691_ ) );
NAND3_X1 \mreg/_08597_ ( .A1(\mreg/_02485_ ), .A2(\mreg/_03999_ ), .A3(\mreg/_02691_ ), .ZN(\mreg/_02692_ ) );
AND4_X1 \mreg/_08598_ ( .A1(\mreg/_02687_ ), .A2(\mreg/_02689_ ), .A3(\mreg/_02690_ ), .A4(\mreg/_02692_ ), .ZN(\mreg/_02693_ ) );
NAND3_X1 \mreg/_08599_ ( .A1(\mreg/_02479_ ), .A2(\mreg/_04031_ ), .A3(\mreg/_02664_ ), .ZN(\mreg/_02694_ ) );
NAND3_X1 \mreg/_08600_ ( .A1(\mreg/_02431_ ), .A2(\mreg/_04095_ ), .A3(\mreg/_02633_ ), .ZN(\mreg/_02695_ ) );
BUF_X4 \mreg/_08601_ ( .A(\mreg/_02597_ ), .Z(\mreg/_02696_ ) );
BUF_X2 \mreg/_08602_ ( .A(\mreg/_02411_ ), .Z(\mreg/_02697_ ) );
NAND3_X1 \mreg/_08603_ ( .A1(\mreg/_02696_ ), .A2(\mreg/_04063_ ), .A3(\mreg/_02697_ ), .ZN(\mreg/_02698_ ) );
BUF_X4 \mreg/_08604_ ( .A(\mreg/_02424_ ), .Z(\mreg/_02699_ ) );
BUF_X2 \mreg/_08605_ ( .A(\mreg/_02553_ ), .Z(\mreg/_02700_ ) );
NAND3_X1 \mreg/_08606_ ( .A1(\mreg/_02699_ ), .A2(\mreg/_04127_ ), .A3(\mreg/_02700_ ), .ZN(\mreg/_02701_ ) );
AND4_X1 \mreg/_08607_ ( .A1(\mreg/_02694_ ), .A2(\mreg/_02695_ ), .A3(\mreg/_02698_ ), .A4(\mreg/_02701_ ), .ZN(\mreg/_02702_ ) );
AND4_X1 \mreg/_08608_ ( .A1(\mreg/_02680_ ), .A2(\mreg/_02686_ ), .A3(\mreg/_02693_ ), .A4(\mreg/_02702_ ), .ZN(\mreg/_02703_ ) );
NAND4_X1 \mreg/_08609_ ( .A1(\mreg/_02667_ ), .A2(\mreg/_02671_ ), .A3(\mreg/_02678_ ), .A4(\mreg/_02703_ ), .ZN(\mreg/_03903_ ) );
NAND3_X1 \mreg/_08610_ ( .A1(\mreg/_02530_ ), .A2(\mreg/_04576_ ), .A3(\mreg/_02532_ ), .ZN(\mreg/_02704_ ) );
NAND3_X1 \mreg/_08611_ ( .A1(\mreg/_02432_ ), .A2(\mreg/_04672_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02705_ ) );
NAND3_X1 \mreg/_08612_ ( .A1(\mreg/_02441_ ), .A2(\mreg/_04608_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02706_ ) );
NAND3_X1 \mreg/_08613_ ( .A1(\mreg/_02426_ ), .A2(\mreg/_01370_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02707_ ) );
AND4_X1 \mreg/_08614_ ( .A1(\mreg/_02704_ ), .A2(\mreg/_02705_ ), .A3(\mreg/_02706_ ), .A4(\mreg/_02707_ ), .ZN(\mreg/_02708_ ) );
NAND4_X1 \mreg/_08615_ ( .A1(\mreg/_02535_ ), .A2(\mreg/_02536_ ), .A3(\mreg/_04512_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_02709_ ) );
OAI21_X1 \mreg/_08616_ ( .A(\mreg/_02709_ ), .B1(\mreg/_02660_ ), .B2(\mreg/_01368_ ), .ZN(\mreg/_02710_ ) );
AOI221_X4 \mreg/_08617_ ( .A(\mreg/_02710_ ), .B1(\mreg/_04480_ ), .B2(\mreg/_02542_ ), .C1(\mreg/_04448_ ), .C2(\mreg/_02544_ ), .ZN(\mreg/_02711_ ) );
NAND4_X1 \mreg/_08618_ ( .A1(\mreg/_02608_ ), .A2(\mreg/_04224_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02609_ ), .ZN(\mreg/_02712_ ) );
OAI21_X1 \mreg/_08619_ ( .A(\mreg/_02712_ ), .B1(\mreg/_02611_ ), .B2(\mreg/_01375_ ), .ZN(\mreg/_02713_ ) );
AOI221_X4 \mreg/_08620_ ( .A(\mreg/_02713_ ), .B1(\mreg/_04192_ ), .B2(\mreg/_02613_ ), .C1(\mreg/_04160_ ), .C2(\mreg/_02614_ ), .ZN(\mreg/_02714_ ) );
BUF_X4 \mreg/_08621_ ( .A(\mreg/_02454_ ), .Z(\mreg/_02715_ ) );
NAND3_X1 \mreg/_08622_ ( .A1(\mreg/_02715_ ), .A2(\mreg/_04384_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02716_ ) );
NAND3_X1 \mreg/_08623_ ( .A1(\mreg/_02459_ ), .A2(\mreg/_04416_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02717_ ) );
NAND3_X1 \mreg/_08624_ ( .A1(\mreg/_02463_ ), .A2(\mreg/_04352_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02718_ ) );
NAND3_X1 \mreg/_08625_ ( .A1(\mreg/_02619_ ), .A2(\mreg/_04320_ ), .A3(\mreg/_02467_ ), .ZN(\mreg/_02719_ ) );
AND4_X1 \mreg/_08626_ ( .A1(\mreg/_02716_ ), .A2(\mreg/_02717_ ), .A3(\mreg/_02718_ ), .A4(\mreg/_02719_ ), .ZN(\mreg/_02720_ ) );
AND4_X4 \mreg/_08627_ ( .A1(\mreg/_02708_ ), .A2(\mreg/_02711_ ), .A3(\mreg/_02714_ ), .A4(\mreg/_02720_ ), .ZN(\mreg/_02721_ ) );
AND3_X1 \mreg/_08628_ ( .A1(\mreg/_02419_ ), .A2(\mreg/_04288_ ), .A3(\mreg/_02697_ ), .ZN(\mreg/_02722_ ) );
BUF_X4 \mreg/_08629_ ( .A(\mreg/_02416_ ), .Z(\mreg/_02723_ ) );
BUF_X4 \mreg/_08630_ ( .A(\mreg/_02627_ ), .Z(\mreg/_02724_ ) );
AOI221_X4 \mreg/_08631_ ( .A(\mreg/_02722_ ), .B1(\mreg/_02723_ ), .B2(\mreg/_04736_ ), .C1(\mreg/_04640_ ), .C2(\mreg/_02724_ ), .ZN(\mreg/_02725_ ) );
NAND3_X1 \mreg/_08632_ ( .A1(\mreg/_02504_ ), .A2(\mreg/_04800_ ), .A3(\mreg/_02624_ ), .ZN(\mreg/_02726_ ) );
NAND3_X1 \mreg/_08633_ ( .A1(\mreg/_02506_ ), .A2(\mreg/_04832_ ), .A3(\mreg/_02642_ ), .ZN(\mreg/_02727_ ) );
NAND3_X1 \mreg/_08634_ ( .A1(\mreg/_02508_ ), .A2(\mreg/_04864_ ), .A3(\mreg/_02652_ ), .ZN(\mreg/_02728_ ) );
BUF_X2 \mreg/_08635_ ( .A(\mreg/_02443_ ), .Z(\mreg/_02729_ ) );
BUF_X2 \mreg/_08636_ ( .A(\mreg/_02729_ ), .Z(\mreg/_02730_ ) );
NAND3_X1 \mreg/_08637_ ( .A1(\mreg/_02730_ ), .A2(\mreg/_02513_ ), .A3(\mreg/_04768_ ), .ZN(\mreg/_02731_ ) );
AND4_X1 \mreg/_08638_ ( .A1(\mreg/_02726_ ), .A2(\mreg/_02727_ ), .A3(\mreg/_02728_ ), .A4(\mreg/_02731_ ), .ZN(\mreg/_02732_ ) );
AND3_X1 \mreg/_08639_ ( .A1(\mreg/_02444_ ), .A2(\mreg/_04896_ ), .A3(\mreg/_02480_ ), .ZN(\mreg/_02733_ ) );
AND2_X1 \mreg/_08640_ ( .A1(\mreg/_02470_ ), .A2(\mreg/_02415_ ), .ZN(\mreg/_02734_ ) );
BUF_X4 \mreg/_08641_ ( .A(\mreg/_02734_ ), .Z(\mreg/_02735_ ) );
AOI21_X1 \mreg/_08642_ ( .A(\mreg/_02733_ ), .B1(\mreg/_02735_ ), .B2(\mreg/_04928_ ), .ZN(\mreg/_02736_ ) );
BUF_X2 \mreg/_08643_ ( .A(\mreg/_02427_ ), .Z(\mreg/_02737_ ) );
NAND3_X1 \mreg/_08644_ ( .A1(\mreg/_02477_ ), .A2(\mreg/_03968_ ), .A3(\mreg/_02737_ ), .ZN(\mreg/_02738_ ) );
NAND2_X4 \mreg/_08645_ ( .A1(\mreg/_02484_ ), .A2(\mreg/_02410_ ), .ZN(\mreg/_02739_ ) );
OAI211_X2 \mreg/_08646_ ( .A(\mreg/_02736_ ), .B(\mreg/_02738_ ), .C1(\mreg/_01395_ ), .C2(\mreg/_02739_ ), .ZN(\mreg/_02740_ ) );
BUF_X2 \mreg/_08647_ ( .A(\mreg/_02444_ ), .Z(\mreg/_02741_ ) );
BUF_X2 \mreg/_08648_ ( .A(\mreg/_02447_ ), .Z(\mreg/_02742_ ) );
AND3_X1 \mreg/_08649_ ( .A1(\mreg/_02741_ ), .A2(\mreg/_04032_ ), .A3(\mreg/_02742_ ), .ZN(\mreg/_02743_ ) );
BUF_X2 \mreg/_08650_ ( .A(\mreg/_02440_ ), .Z(\mreg/_02744_ ) );
CLKBUF_X2 \mreg/_08651_ ( .A(\mreg/_02427_ ), .Z(\mreg/_02745_ ) );
AND3_X1 \mreg/_08652_ ( .A1(\mreg/_02744_ ), .A2(\mreg/_04064_ ), .A3(\mreg/_02745_ ), .ZN(\mreg/_02746_ ) );
BUF_X4 \mreg/_08653_ ( .A(\mreg/_02427_ ), .Z(\mreg/_02747_ ) );
NAND3_X1 \mreg/_08654_ ( .A1(\mreg/_02426_ ), .A2(\mreg/_04128_ ), .A3(\mreg/_02747_ ), .ZN(\mreg/_02748_ ) );
NAND2_X1 \mreg/_08655_ ( .A1(\mreg/_02430_ ), .A2(\mreg/_02410_ ), .ZN(\mreg/_02749_ ) );
OAI21_X1 \mreg/_08656_ ( .A(\mreg/_02748_ ), .B1(\mreg/_02749_ ), .B2(\mreg/_01394_ ), .ZN(\mreg/_02750_ ) );
NOR4_X1 \mreg/_08657_ ( .A1(\mreg/_02740_ ), .A2(\mreg/_02743_ ), .A3(\mreg/_02746_ ), .A4(\mreg/_02750_ ), .ZN(\mreg/_02751_ ) );
NAND4_X1 \mreg/_08658_ ( .A1(\mreg/_02721_ ), .A2(\mreg/_02725_ ), .A3(\mreg/_02732_ ), .A4(\mreg/_02751_ ), .ZN(\mreg/_03904_ ) );
NAND3_X1 \mreg/_08659_ ( .A1(\mreg/_02530_ ), .A2(\mreg/_04577_ ), .A3(\mreg/_02532_ ), .ZN(\mreg/_02752_ ) );
NAND3_X1 \mreg/_08660_ ( .A1(\mreg/_02432_ ), .A2(\mreg/_04673_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02753_ ) );
NAND3_X1 \mreg/_08661_ ( .A1(\mreg/_02441_ ), .A2(\mreg/_04609_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02754_ ) );
NAND3_X1 \mreg/_08662_ ( .A1(\mreg/_02426_ ), .A2(\mreg/_01416_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02755_ ) );
AND4_X1 \mreg/_08663_ ( .A1(\mreg/_02752_ ), .A2(\mreg/_02753_ ), .A3(\mreg/_02754_ ), .A4(\mreg/_02755_ ), .ZN(\mreg/_02756_ ) );
NAND4_X1 \mreg/_08664_ ( .A1(\mreg/_02535_ ), .A2(\mreg/_02536_ ), .A3(\mreg/_04513_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_02757_ ) );
OAI21_X1 \mreg/_08665_ ( .A(\mreg/_02757_ ), .B1(\mreg/_02660_ ), .B2(\mreg/_01410_ ), .ZN(\mreg/_02758_ ) );
BUF_X4 \mreg/_08666_ ( .A(\mreg/_02541_ ), .Z(\mreg/_02759_ ) );
BUF_X4 \mreg/_08667_ ( .A(\mreg/_02543_ ), .Z(\mreg/_02760_ ) );
AOI221_X4 \mreg/_08668_ ( .A(\mreg/_02758_ ), .B1(\mreg/_04481_ ), .B2(\mreg/_02759_ ), .C1(\mreg/_04449_ ), .C2(\mreg/_02760_ ), .ZN(\mreg/_02761_ ) );
NAND4_X1 \mreg/_08669_ ( .A1(\mreg/_02608_ ), .A2(\mreg/_04225_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02609_ ), .ZN(\mreg/_02762_ ) );
OAI21_X1 \mreg/_08670_ ( .A(\mreg/_02762_ ), .B1(\mreg/_02611_ ), .B2(\mreg/_01421_ ), .ZN(\mreg/_02763_ ) );
AOI221_X4 \mreg/_08671_ ( .A(\mreg/_02763_ ), .B1(\mreg/_04193_ ), .B2(\mreg/_02613_ ), .C1(\mreg/_04161_ ), .C2(\mreg/_02614_ ), .ZN(\mreg/_02764_ ) );
NAND3_X1 \mreg/_08672_ ( .A1(\mreg/_02715_ ), .A2(\mreg/_04385_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02765_ ) );
NAND3_X1 \mreg/_08673_ ( .A1(\mreg/_02565_ ), .A2(\mreg/_04417_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02766_ ) );
BUF_X2 \mreg/_08674_ ( .A(\mreg/_02462_ ), .Z(\mreg/_02767_ ) );
NAND3_X1 \mreg/_08675_ ( .A1(\mreg/_02767_ ), .A2(\mreg/_04353_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02768_ ) );
NAND3_X1 \mreg/_08676_ ( .A1(\mreg/_02619_ ), .A2(\mreg/_04321_ ), .A3(\mreg/_02467_ ), .ZN(\mreg/_02769_ ) );
AND4_X1 \mreg/_08677_ ( .A1(\mreg/_02765_ ), .A2(\mreg/_02766_ ), .A3(\mreg/_02768_ ), .A4(\mreg/_02769_ ), .ZN(\mreg/_02770_ ) );
AND4_X4 \mreg/_08678_ ( .A1(\mreg/_02756_ ), .A2(\mreg/_02761_ ), .A3(\mreg/_02764_ ), .A4(\mreg/_02770_ ), .ZN(\mreg/_02771_ ) );
AND3_X1 \mreg/_08679_ ( .A1(\mreg/_02419_ ), .A2(\mreg/_04289_ ), .A3(\mreg/_02697_ ), .ZN(\mreg/_02772_ ) );
AOI221_X4 \mreg/_08680_ ( .A(\mreg/_02772_ ), .B1(\mreg/_02723_ ), .B2(\mreg/_04737_ ), .C1(\mreg/_04641_ ), .C2(\mreg/_02724_ ), .ZN(\mreg/_02773_ ) );
NAND3_X1 \mreg/_08681_ ( .A1(\mreg/_02504_ ), .A2(\mreg/_04801_ ), .A3(\mreg/_02624_ ), .ZN(\mreg/_02774_ ) );
NAND3_X1 \mreg/_08682_ ( .A1(\mreg/_02506_ ), .A2(\mreg/_04833_ ), .A3(\mreg/_02642_ ), .ZN(\mreg/_02775_ ) );
NAND3_X1 \mreg/_08683_ ( .A1(\mreg/_02508_ ), .A2(\mreg/_04865_ ), .A3(\mreg/_02652_ ), .ZN(\mreg/_02776_ ) );
NAND3_X1 \mreg/_08684_ ( .A1(\mreg/_02730_ ), .A2(\mreg/_02513_ ), .A3(\mreg/_04769_ ), .ZN(\mreg/_02777_ ) );
AND4_X1 \mreg/_08685_ ( .A1(\mreg/_02774_ ), .A2(\mreg/_02775_ ), .A3(\mreg/_02776_ ), .A4(\mreg/_02777_ ), .ZN(\mreg/_02778_ ) );
BUF_X4 \mreg/_08686_ ( .A(\mreg/_02434_ ), .Z(\mreg/_02779_ ) );
NAND3_X1 \mreg/_08687_ ( .A1(\mreg/_02477_ ), .A2(\mreg/_03969_ ), .A3(\mreg/_02779_ ), .ZN(\mreg/_02780_ ) );
NAND3_X1 \mreg/_08688_ ( .A1(\mreg/_02647_ ), .A2(\mreg/_04001_ ), .A3(\mreg/_02737_ ), .ZN(\mreg/_02781_ ) );
NAND3_X1 \mreg/_08689_ ( .A1(\mreg/_02472_ ), .A2(\mreg/_04929_ ), .A3(\mreg/_02737_ ), .ZN(\mreg/_02782_ ) );
NAND3_X1 \mreg/_08690_ ( .A1(\mreg/_02741_ ), .A2(\mreg/_02645_ ), .A3(\mreg/_04897_ ), .ZN(\mreg/_02783_ ) );
NAND4_X1 \mreg/_08691_ ( .A1(\mreg/_02780_ ), .A2(\mreg/_02781_ ), .A3(\mreg/_02782_ ), .A4(\mreg/_02783_ ), .ZN(\mreg/_02784_ ) );
BUF_X2 \mreg/_08692_ ( .A(\mreg/_02431_ ), .Z(\mreg/_02785_ ) );
NAND3_X1 \mreg/_08693_ ( .A1(\mreg/_02785_ ), .A2(\mreg/_04097_ ), .A3(\mreg/_02737_ ), .ZN(\mreg/_02786_ ) );
BUF_X2 \mreg/_08694_ ( .A(\mreg/_02425_ ), .Z(\mreg/_02787_ ) );
NAND3_X1 \mreg/_08695_ ( .A1(\mreg/_02787_ ), .A2(\mreg/_04129_ ), .A3(\mreg/_02737_ ), .ZN(\mreg/_02788_ ) );
NAND2_X1 \mreg/_08696_ ( .A1(\mreg/_02786_ ), .A2(\mreg/_02788_ ), .ZN(\mreg/_02789_ ) );
AND3_X1 \mreg/_08697_ ( .A1(\mreg/_02741_ ), .A2(\mreg/_04033_ ), .A3(\mreg/_02532_ ), .ZN(\mreg/_02790_ ) );
AND3_X1 \mreg/_08698_ ( .A1(\mreg/_02744_ ), .A2(\mreg/_04065_ ), .A3(\mreg/_02745_ ), .ZN(\mreg/_02791_ ) );
NOR4_X1 \mreg/_08699_ ( .A1(\mreg/_02784_ ), .A2(\mreg/_02789_ ), .A3(\mreg/_02790_ ), .A4(\mreg/_02791_ ), .ZN(\mreg/_02792_ ) );
NAND4_X1 \mreg/_08700_ ( .A1(\mreg/_02771_ ), .A2(\mreg/_02773_ ), .A3(\mreg/_02778_ ), .A4(\mreg/_02792_ ), .ZN(\mreg/_03905_ ) );
NAND3_X1 \mreg/_08701_ ( .A1(\mreg/_02531_ ), .A2(\mreg/_04578_ ), .A3(\mreg/_02533_ ), .ZN(\mreg/_02793_ ) );
NAND4_X1 \mreg/_08702_ ( .A1(\mreg/_02535_ ), .A2(\mreg/_02536_ ), .A3(\mreg/_04514_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_02794_ ) );
OAI21_X1 \mreg/_08703_ ( .A(\mreg/_02794_ ), .B1(\mreg/_02660_ ), .B2(\mreg/_01455_ ), .ZN(\mreg/_02795_ ) );
AOI221_X4 \mreg/_08704_ ( .A(\mreg/_02795_ ), .B1(\mreg/_04482_ ), .B2(\mreg/_02759_ ), .C1(\mreg/_04450_ ), .C2(\mreg/_02760_ ), .ZN(\mreg/_02796_ ) );
NAND3_X1 \mreg/_08705_ ( .A1(\mreg/_02546_ ), .A2(\mreg/_04610_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02797_ ) );
AND3_X1 \mreg/_08706_ ( .A1(\mreg/_02432_ ), .A2(\mreg/_04674_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02798_ ) );
AOI21_X1 \mreg/_08707_ ( .A(\mreg/_02798_ ), .B1(\mreg/_01450_ ), .B2(\mreg/_02550_ ), .ZN(\mreg/_02799_ ) );
AND4_X4 \mreg/_08708_ ( .A1(\mreg/_02793_ ), .A2(\mreg/_02796_ ), .A3(\mreg/_02797_ ), .A4(\mreg/_02799_ ), .ZN(\mreg/_02800_ ) );
NAND3_X1 \mreg/_08709_ ( .A1(\mreg/_02672_ ), .A2(\mreg/_04386_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02801_ ) );
NAND4_X1 \mreg/_08710_ ( .A1(\mreg/_02608_ ), .A2(\mreg/_04226_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02499_ ), .ZN(\mreg/_02802_ ) );
OAI21_X1 \mreg/_08711_ ( .A(\mreg/_02802_ ), .B1(\mreg/_02611_ ), .B2(\mreg/_01463_ ), .ZN(\mreg/_02803_ ) );
AOI221_X4 \mreg/_08712_ ( .A(\mreg/_02803_ ), .B1(\mreg/_04194_ ), .B2(\mreg/_02613_ ), .C1(\mreg/_04162_ ), .C2(\mreg/_02614_ ), .ZN(\mreg/_02804_ ) );
NAND3_X1 \mreg/_08713_ ( .A1(\mreg/_02674_ ), .A2(\mreg/_04418_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02805_ ) );
AND3_X1 \mreg/_08714_ ( .A1(\mreg/_02767_ ), .A2(\mreg/_04354_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02806_ ) );
AND2_X2 \mreg/_08715_ ( .A1(\mreg/_02510_ ), .A2(\mreg/_02466_ ), .ZN(\mreg/_02807_ ) );
AOI21_X1 \mreg/_08716_ ( .A(\mreg/_02806_ ), .B1(\mreg/_04322_ ), .B2(\mreg/_02807_ ), .ZN(\mreg/_02808_ ) );
AND4_X1 \mreg/_08717_ ( .A1(\mreg/_02801_ ), .A2(\mreg/_02804_ ), .A3(\mreg/_02805_ ), .A4(\mreg/_02808_ ), .ZN(\mreg/_02809_ ) );
NAND3_X1 \mreg/_08718_ ( .A1(\mreg/_02583_ ), .A2(\mreg/_04290_ ), .A3(\mreg/_02624_ ), .ZN(\mreg/_02810_ ) );
AND3_X1 \mreg/_08719_ ( .A1(\mreg/_02565_ ), .A2(\mreg/_04866_ ), .A3(\mreg/_02566_ ), .ZN(\mreg/_02811_ ) );
AOI21_X1 \mreg/_08720_ ( .A(\mreg/_02811_ ), .B1(\mreg/_04834_ ), .B2(\mreg/_02636_ ), .ZN(\mreg/_02812_ ) );
AOI22_X1 \mreg/_08721_ ( .A1(\mreg/_04642_ ), .A2(\mreg/_02724_ ), .B1(\mreg/_02723_ ), .B2(\mreg/_04738_ ), .ZN(\mreg/_02813_ ) );
AND2_X2 \mreg/_08722_ ( .A1(\mreg/_02462_ ), .A2(\mreg/_02410_ ), .ZN(\mreg/_02814_ ) );
BUF_X4 \mreg/_08723_ ( .A(\mreg/_02814_ ), .Z(\mreg/_02815_ ) );
AND2_X1 \mreg/_08724_ ( .A1(\mreg/_02443_ ), .A2(\mreg/_02452_ ), .ZN(\mreg/_02816_ ) );
BUF_X4 \mreg/_08725_ ( .A(\mreg/_02816_ ), .Z(\mreg/_02817_ ) );
AOI22_X1 \mreg/_08726_ ( .A1(\mreg/_02815_ ), .A2(\mreg/_04802_ ), .B1(\mreg/_04770_ ), .B2(\mreg/_02817_ ), .ZN(\mreg/_02818_ ) );
AND4_X1 \mreg/_08727_ ( .A1(\mreg/_02810_ ), .A2(\mreg/_02812_ ), .A3(\mreg/_02813_ ), .A4(\mreg/_02818_ ), .ZN(\mreg/_02819_ ) );
BUF_X4 \mreg/_08728_ ( .A(\mreg/_02623_ ), .Z(\mreg/_02820_ ) );
NAND3_X1 \mreg/_08729_ ( .A1(\mreg/_02641_ ), .A2(\mreg/_03970_ ), .A3(\mreg/_02820_ ), .ZN(\mreg/_02821_ ) );
NAND3_X1 \mreg/_08730_ ( .A1(\mreg/_02629_ ), .A2(\mreg/_04034_ ), .A3(\mreg/_02448_ ), .ZN(\mreg/_02822_ ) );
NAND3_X1 \mreg/_08731_ ( .A1(\mreg/_02571_ ), .A2(\mreg/_04098_ ), .A3(\mreg/_02486_ ), .ZN(\mreg/_02823_ ) );
NAND3_X1 \mreg/_08732_ ( .A1(\mreg/_02696_ ), .A2(\mreg/_04066_ ), .A3(\mreg/_02572_ ), .ZN(\mreg/_02824_ ) );
NAND3_X1 \mreg/_08733_ ( .A1(\mreg/_02699_ ), .A2(\mreg/_04130_ ), .A3(\mreg/_02633_ ), .ZN(\mreg/_02825_ ) );
AND4_X1 \mreg/_08734_ ( .A1(\mreg/_02822_ ), .A2(\mreg/_02823_ ), .A3(\mreg/_02824_ ), .A4(\mreg/_02825_ ), .ZN(\mreg/_02826_ ) );
NAND3_X1 \mreg/_08735_ ( .A1(\mreg/_02647_ ), .A2(\mreg/_04002_ ), .A3(\mreg/_02654_ ), .ZN(\mreg/_02827_ ) );
AND3_X1 \mreg/_08736_ ( .A1(\mreg/_02729_ ), .A2(\mreg/_04898_ ), .A3(\mreg/_02644_ ), .ZN(\mreg/_02828_ ) );
AOI21_X1 \mreg/_08737_ ( .A(\mreg/_02828_ ), .B1(\mreg/_02735_ ), .B2(\mreg/_04930_ ), .ZN(\mreg/_02829_ ) );
AND4_X1 \mreg/_08738_ ( .A1(\mreg/_02821_ ), .A2(\mreg/_02826_ ), .A3(\mreg/_02827_ ), .A4(\mreg/_02829_ ), .ZN(\mreg/_02830_ ) );
NAND4_X1 \mreg/_08739_ ( .A1(\mreg/_02800_ ), .A2(\mreg/_02809_ ), .A3(\mreg/_02819_ ), .A4(\mreg/_02830_ ), .ZN(\mreg/_03906_ ) );
NAND3_X1 \mreg/_08740_ ( .A1(\mreg/_02785_ ), .A2(\mreg/_04099_ ), .A3(\mreg/_02779_ ), .ZN(\mreg/_02831_ ) );
NAND3_X1 \mreg/_08741_ ( .A1(\mreg/_02730_ ), .A2(\mreg/_04035_ ), .A3(\mreg/_02742_ ), .ZN(\mreg/_02832_ ) );
OAI211_X2 \mreg/_08742_ ( .A(\mreg/_02831_ ), .B(\mreg/_02832_ ), .C1(\mreg/_02739_ ), .C2(\mreg/_01516_ ), .ZN(\mreg/_02833_ ) );
NAND3_X1 \mreg/_08743_ ( .A1(\mreg/_02639_ ), .A2(\mreg/_04483_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02834_ ) );
NAND3_X1 \mreg/_08744_ ( .A1(\mreg/_02744_ ), .A2(\mreg/_04611_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02835_ ) );
NAND3_X1 \mreg/_08745_ ( .A1(\mreg/_02511_ ), .A2(\mreg/_04579_ ), .A3(\mreg/_02532_ ), .ZN(\mreg/_02836_ ) );
BUF_X2 \mreg/_08746_ ( .A(\mreg/_02510_ ), .Z(\mreg/_02837_ ) );
BUF_X2 \mreg/_08747_ ( .A(\mreg/_02480_ ), .Z(\mreg/_02838_ ) );
NAND3_X1 \mreg/_08748_ ( .A1(\mreg/_02837_ ), .A2(\mreg/_04451_ ), .A3(\mreg/_02838_ ), .ZN(\mreg/_02839_ ) );
NAND4_X1 \mreg/_08749_ ( .A1(\mreg/_02834_ ), .A2(\mreg/_02835_ ), .A3(\mreg/_02836_ ), .A4(\mreg/_02839_ ), .ZN(\mreg/_02840_ ) );
NAND3_X1 \mreg/_08750_ ( .A1(\mreg/_02455_ ), .A2(\mreg/_04387_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02841_ ) );
BUF_X2 \mreg/_08751_ ( .A(\mreg/_02458_ ), .Z(\mreg/_02842_ ) );
NAND3_X1 \mreg/_08752_ ( .A1(\mreg/_02842_ ), .A2(\mreg/_04419_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02843_ ) );
NAND3_X1 \mreg/_08753_ ( .A1(\mreg/_02837_ ), .A2(\mreg/_04163_ ), .A3(\mreg/_02581_ ), .ZN(\mreg/_02844_ ) );
BUF_X2 \mreg/_08754_ ( .A(\mreg/_02419_ ), .Z(\mreg/_02845_ ) );
NAND3_X1 \mreg/_08755_ ( .A1(\mreg/_02845_ ), .A2(\mreg/_04195_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02846_ ) );
NAND4_X1 \mreg/_08756_ ( .A1(\mreg/_02841_ ), .A2(\mreg/_02843_ ), .A3(\mreg/_02844_ ), .A4(\mreg/_02846_ ), .ZN(\mreg/_02847_ ) );
NAND3_X1 \mreg/_08757_ ( .A1(\mreg/_02842_ ), .A2(\mreg/_04867_ ), .A3(\mreg/_02745_ ), .ZN(\mreg/_02848_ ) );
NAND3_X1 \mreg/_08758_ ( .A1(\mreg/_02845_ ), .A2(\mreg/_04291_ ), .A3(\mreg/_02745_ ), .ZN(\mreg/_02849_ ) );
NAND3_X1 \mreg/_08759_ ( .A1(\mreg/_02490_ ), .A2(\mreg/_04643_ ), .A3(\mreg/_02747_ ), .ZN(\mreg/_02850_ ) );
BUF_X2 \mreg/_08760_ ( .A(\mreg/_02480_ ), .Z(\mreg/_02851_ ) );
NAND3_X1 \mreg/_08761_ ( .A1(\mreg/_02741_ ), .A2(\mreg/_02851_ ), .A3(\mreg/_04899_ ), .ZN(\mreg/_02852_ ) );
NAND4_X1 \mreg/_08762_ ( .A1(\mreg/_02848_ ), .A2(\mreg/_02849_ ), .A3(\mreg/_02850_ ), .A4(\mreg/_02852_ ), .ZN(\mreg/_02853_ ) );
NOR4_X1 \mreg/_08763_ ( .A1(\mreg/_02833_ ), .A2(\mreg/_02840_ ), .A3(\mreg/_02847_ ), .A4(\mreg/_02853_ ), .ZN(\mreg/_02854_ ) );
CLKBUF_X2 \mreg/_08764_ ( .A(\mreg/_02414_ ), .Z(\mreg/_02855_ ) );
NAND3_X1 \mreg/_08765_ ( .A1(\mreg/_02855_ ), .A2(\mreg/_04739_ ), .A3(\mreg/_02633_ ), .ZN(\mreg/_02856_ ) );
NAND3_X1 \mreg/_08766_ ( .A1(\mreg/_02729_ ), .A2(\mreg/_02466_ ), .A3(\mreg/_04771_ ), .ZN(\mreg/_02857_ ) );
NAND2_X1 \mreg/_08767_ ( .A1(\mreg/_02856_ ), .A2(\mreg/_02857_ ), .ZN(\mreg/_02858_ ) );
AOI221_X4 \mreg/_08768_ ( .A(\mreg/_02858_ ), .B1(\mreg/_04803_ ), .B2(\mreg/_02814_ ), .C1(\mreg/_04835_ ), .C2(\mreg/_02636_ ), .ZN(\mreg/_02859_ ) );
NAND3_X1 \mreg/_08769_ ( .A1(\mreg/_02785_ ), .A2(\mreg/_04675_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02860_ ) );
NAND3_X1 \mreg/_08770_ ( .A1(\mreg/_02787_ ), .A2(\mreg/_01488_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02861_ ) );
NAND4_X1 \mreg/_08771_ ( .A1(\mreg/_02587_ ), .A2(\mreg/_02838_ ), .A3(\mreg/_04515_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_02862_ ) );
NAND4_X1 \mreg/_08772_ ( .A1(\mreg/_02645_ ), .A2(\mreg/_04547_ ), .A3(\mreg/_02589_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_02863_ ) );
NAND4_X1 \mreg/_08773_ ( .A1(\mreg/_02860_ ), .A2(\mreg/_02861_ ), .A3(\mreg/_02862_ ), .A4(\mreg/_02863_ ), .ZN(\mreg/_02864_ ) );
NAND4_X1 \mreg/_08774_ ( .A1(\mreg/_02587_ ), .A2(\mreg/_04227_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02581_ ), .ZN(\mreg/_02865_ ) );
OAI21_X1 \mreg/_08775_ ( .A(\mreg/_02865_ ), .B1(\mreg/_02493_ ), .B2(\mreg/_01503_ ), .ZN(\mreg/_02866_ ) );
AND3_X1 \mreg/_08776_ ( .A1(\mreg/_02503_ ), .A2(\mreg/_04355_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02867_ ) );
AND3_X1 \mreg/_08777_ ( .A1(\mreg/_02837_ ), .A2(\mreg/_04323_ ), .A3(\mreg/_02512_ ), .ZN(\mreg/_02868_ ) );
NOR4_X1 \mreg/_08778_ ( .A1(\mreg/_02864_ ), .A2(\mreg/_02866_ ), .A3(\mreg/_02867_ ), .A4(\mreg/_02868_ ), .ZN(\mreg/_02869_ ) );
NAND3_X1 \mreg/_08779_ ( .A1(\mreg/_02639_ ), .A2(\mreg/_04931_ ), .A3(\mreg/_02820_ ), .ZN(\mreg/_02870_ ) );
NAND3_X1 \mreg/_08780_ ( .A1(\mreg/_02641_ ), .A2(\mreg/_03971_ ), .A3(\mreg/_02652_ ), .ZN(\mreg/_02871_ ) );
NAND3_X1 \mreg/_08781_ ( .A1(\mreg/_02744_ ), .A2(\mreg/_04067_ ), .A3(\mreg/_02654_ ), .ZN(\mreg/_02872_ ) );
NAND3_X1 \mreg/_08782_ ( .A1(\mreg/_02787_ ), .A2(\mreg/_04131_ ), .A3(\mreg/_02648_ ), .ZN(\mreg/_02873_ ) );
AND4_X1 \mreg/_08783_ ( .A1(\mreg/_02870_ ), .A2(\mreg/_02871_ ), .A3(\mreg/_02872_ ), .A4(\mreg/_02873_ ), .ZN(\mreg/_02874_ ) );
NAND4_X1 \mreg/_08784_ ( .A1(\mreg/_02854_ ), .A2(\mreg/_02859_ ), .A3(\mreg/_02869_ ), .A4(\mreg/_02874_ ), .ZN(\mreg/_03907_ ) );
NAND3_X1 \mreg/_08785_ ( .A1(\mreg/_02597_ ), .A2(\mreg/_04612_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02875_ ) );
NAND3_X1 \mreg/_08786_ ( .A1(\mreg/_02599_ ), .A2(\mreg/_04580_ ), .A3(\mreg/_02446_ ), .ZN(\mreg/_02876_ ) );
NAND2_X1 \mreg/_08787_ ( .A1(\mreg/_02875_ ), .A2(\mreg/_02876_ ), .ZN(\mreg/_02877_ ) );
AOI221_X4 \mreg/_08788_ ( .A(\mreg/_02877_ ), .B1(\mreg/_01531_ ), .B2(\mreg/_02549_ ), .C1(\mreg/_04676_ ), .C2(\mreg/_02603_ ), .ZN(\mreg/_02878_ ) );
BUF_X4 \mreg/_08789_ ( .A(\mreg/_02474_ ), .Z(\mreg/_02879_ ) );
NAND4_X1 \mreg/_08790_ ( .A1(\mreg/_02535_ ), .A2(\mreg/_02879_ ), .A3(\mreg/_04516_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_02880_ ) );
OAI21_X1 \mreg/_08791_ ( .A(\mreg/_02880_ ), .B1(\mreg/_02660_ ), .B2(\mreg/_01529_ ), .ZN(\mreg/_02881_ ) );
AOI221_X4 \mreg/_08792_ ( .A(\mreg/_02881_ ), .B1(\mreg/_04484_ ), .B2(\mreg/_02759_ ), .C1(\mreg/_04452_ ), .C2(\mreg/_02760_ ), .ZN(\mreg/_02882_ ) );
NAND4_X1 \mreg/_08793_ ( .A1(\mreg/_02608_ ), .A2(\mreg/_04228_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02499_ ), .ZN(\mreg/_02883_ ) );
OAI21_X1 \mreg/_08794_ ( .A(\mreg/_02883_ ), .B1(\mreg/_02611_ ), .B2(\mreg/_01538_ ), .ZN(\mreg/_02884_ ) );
AOI221_X4 \mreg/_08795_ ( .A(\mreg/_02884_ ), .B1(\mreg/_04196_ ), .B2(\mreg/_02613_ ), .C1(\mreg/_04164_ ), .C2(\mreg/_02614_ ), .ZN(\mreg/_02885_ ) );
NAND3_X1 \mreg/_08796_ ( .A1(\mreg/_02715_ ), .A2(\mreg/_04388_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02886_ ) );
NAND3_X1 \mreg/_08797_ ( .A1(\mreg/_02565_ ), .A2(\mreg/_04420_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02887_ ) );
NAND3_X1 \mreg/_08798_ ( .A1(\mreg/_02767_ ), .A2(\mreg/_04356_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02888_ ) );
NAND3_X1 \mreg/_08799_ ( .A1(\mreg/_02520_ ), .A2(\mreg/_04324_ ), .A3(\mreg/_02467_ ), .ZN(\mreg/_02889_ ) );
AND4_X1 \mreg/_08800_ ( .A1(\mreg/_02886_ ), .A2(\mreg/_02887_ ), .A3(\mreg/_02888_ ), .A4(\mreg/_02889_ ), .ZN(\mreg/_02890_ ) );
AND4_X4 \mreg/_08801_ ( .A1(\mreg/_02878_ ), .A2(\mreg/_02882_ ), .A3(\mreg/_02885_ ), .A4(\mreg/_02890_ ), .ZN(\mreg/_02891_ ) );
AND3_X1 \mreg/_08802_ ( .A1(\mreg/_02490_ ), .A2(\mreg/_04644_ ), .A3(\mreg/_02700_ ), .ZN(\mreg/_02892_ ) );
AOI221_X4 \mreg/_08803_ ( .A(\mreg/_02892_ ), .B1(\mreg/_02723_ ), .B2(\mreg/_04740_ ), .C1(\mreg/_04292_ ), .C2(\mreg/_02421_ ), .ZN(\mreg/_02893_ ) );
NAND3_X1 \mreg/_08804_ ( .A1(\mreg/_02504_ ), .A2(\mreg/_04804_ ), .A3(\mreg/_02624_ ), .ZN(\mreg/_02894_ ) );
NAND3_X1 \mreg/_08805_ ( .A1(\mreg/_02506_ ), .A2(\mreg/_04836_ ), .A3(\mreg/_02642_ ), .ZN(\mreg/_02895_ ) );
NAND3_X1 \mreg/_08806_ ( .A1(\mreg/_02508_ ), .A2(\mreg/_04868_ ), .A3(\mreg/_02654_ ), .ZN(\mreg/_02896_ ) );
NAND3_X1 \mreg/_08807_ ( .A1(\mreg/_02730_ ), .A2(\mreg/_02513_ ), .A3(\mreg/_04772_ ), .ZN(\mreg/_02897_ ) );
AND4_X1 \mreg/_08808_ ( .A1(\mreg/_02894_ ), .A2(\mreg/_02895_ ), .A3(\mreg/_02896_ ), .A4(\mreg/_02897_ ), .ZN(\mreg/_02898_ ) );
AND3_X1 \mreg/_08809_ ( .A1(\mreg/_02444_ ), .A2(\mreg/_04900_ ), .A3(\mreg/_02480_ ), .ZN(\mreg/_02899_ ) );
AOI21_X1 \mreg/_08810_ ( .A(\mreg/_02899_ ), .B1(\mreg/_02735_ ), .B2(\mreg/_04932_ ), .ZN(\mreg/_02900_ ) );
NAND3_X1 \mreg/_08811_ ( .A1(\mreg/_02477_ ), .A2(\mreg/_03972_ ), .A3(\mreg/_02737_ ), .ZN(\mreg/_02901_ ) );
OAI211_X2 \mreg/_08812_ ( .A(\mreg/_02900_ ), .B(\mreg/_02901_ ), .C1(\mreg/_01544_ ), .C2(\mreg/_02739_ ), .ZN(\mreg/_02902_ ) );
AND3_X1 \mreg/_08813_ ( .A1(\mreg/_02741_ ), .A2(\mreg/_04036_ ), .A3(\mreg/_02742_ ), .ZN(\mreg/_02903_ ) );
AND3_X1 \mreg/_08814_ ( .A1(\mreg/_02744_ ), .A2(\mreg/_04068_ ), .A3(\mreg/_02745_ ), .ZN(\mreg/_02904_ ) );
NAND3_X1 \mreg/_08815_ ( .A1(\mreg/_02426_ ), .A2(\mreg/_04132_ ), .A3(\mreg/_02747_ ), .ZN(\mreg/_02905_ ) );
OAI21_X1 \mreg/_08816_ ( .A(\mreg/_02905_ ), .B1(\mreg/_02749_ ), .B2(\mreg/_01543_ ), .ZN(\mreg/_02906_ ) );
NOR4_X1 \mreg/_08817_ ( .A1(\mreg/_02902_ ), .A2(\mreg/_02903_ ), .A3(\mreg/_02904_ ), .A4(\mreg/_02906_ ), .ZN(\mreg/_02907_ ) );
NAND4_X1 \mreg/_08818_ ( .A1(\mreg/_02891_ ), .A2(\mreg/_02893_ ), .A3(\mreg/_02898_ ), .A4(\mreg/_02907_ ), .ZN(\mreg/_03908_ ) );
NAND3_X1 \mreg/_08819_ ( .A1(\mreg/_02516_ ), .A2(\mreg/_04677_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02908_ ) );
NAND4_X1 \mreg/_08820_ ( .A1(\mreg/_02535_ ), .A2(\mreg/_02879_ ), .A3(\mreg/_04517_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_02909_ ) );
OAI21_X1 \mreg/_08821_ ( .A(\mreg/_02909_ ), .B1(\mreg/_02660_ ), .B2(\mreg/_01570_ ), .ZN(\mreg/_02910_ ) );
AOI221_X1 \mreg/_08822_ ( .A(\mreg/_02910_ ), .B1(\mreg/_04485_ ), .B2(\mreg/_02759_ ), .C1(\mreg/_04453_ ), .C2(\mreg/_02760_ ), .ZN(\mreg/_02911_ ) );
NAND3_X1 \mreg/_08823_ ( .A1(\mreg/_02524_ ), .A2(\mreg/_01572_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02912_ ) );
AND3_X1 \mreg/_08824_ ( .A1(\mreg/_02619_ ), .A2(\mreg/_04581_ ), .A3(\mreg/_02664_ ), .ZN(\mreg/_02913_ ) );
AOI21_X1 \mreg/_08825_ ( .A(\mreg/_02913_ ), .B1(\mreg/_02527_ ), .B2(\mreg/_04613_ ), .ZN(\mreg/_02914_ ) );
AND4_X1 \mreg/_08826_ ( .A1(\mreg/_02908_ ), .A2(\mreg/_02911_ ), .A3(\mreg/_02912_ ), .A4(\mreg/_02914_ ), .ZN(\mreg/_02915_ ) );
AND3_X1 \mreg/_08827_ ( .A1(\mreg/_02409_ ), .A2(\mreg/_04645_ ), .A3(\mreg/_02553_ ), .ZN(\mreg/_02916_ ) );
AOI221_X4 \mreg/_08828_ ( .A(\mreg/_02916_ ), .B1(\mreg/_02416_ ), .B2(\mreg/_04741_ ), .C1(\mreg/_04293_ ), .C2(\mreg/_02421_ ), .ZN(\mreg/_02917_ ) );
NAND3_X1 \mreg/_08829_ ( .A1(\mreg/_02453_ ), .A2(\mreg/_04837_ ), .A3(\mreg/_02553_ ), .ZN(\mreg/_02918_ ) );
NAND3_X1 \mreg/_08830_ ( .A1(\mreg/_02458_ ), .A2(\mreg/_04869_ ), .A3(\mreg/_02553_ ), .ZN(\mreg/_02919_ ) );
NAND2_X1 \mreg/_08831_ ( .A1(\mreg/_02918_ ), .A2(\mreg/_02919_ ), .ZN(\mreg/_02920_ ) );
AOI221_X4 \mreg/_08832_ ( .A(\mreg/_02920_ ), .B1(\mreg/_04805_ ), .B2(\mreg/_02814_ ), .C1(\mreg/_04773_ ), .C2(\mreg/_02817_ ), .ZN(\mreg/_02921_ ) );
NAND3_X1 \mreg/_08833_ ( .A1(\mreg/_02472_ ), .A2(\mreg/_04933_ ), .A3(\mreg/_02434_ ), .ZN(\mreg/_02922_ ) );
NAND3_X1 \mreg/_08834_ ( .A1(\mreg/_02477_ ), .A2(\mreg/_03973_ ), .A3(\mreg/_02563_ ), .ZN(\mreg/_02923_ ) );
NAND3_X1 \mreg/_08835_ ( .A1(\mreg/_02479_ ), .A2(\mreg/_02481_ ), .A3(\mreg/_04901_ ), .ZN(\mreg/_02924_ ) );
NAND3_X1 \mreg/_08836_ ( .A1(\mreg/_02485_ ), .A2(\mreg/_04005_ ), .A3(\mreg/_02688_ ), .ZN(\mreg/_02925_ ) );
AND4_X1 \mreg/_08837_ ( .A1(\mreg/_02922_ ), .A2(\mreg/_02923_ ), .A3(\mreg/_02924_ ), .A4(\mreg/_02925_ ), .ZN(\mreg/_02926_ ) );
NAND3_X1 \mreg/_08838_ ( .A1(\mreg/_02445_ ), .A2(\mreg/_04037_ ), .A3(\mreg/_02448_ ), .ZN(\mreg/_02927_ ) );
NAND3_X1 \mreg/_08839_ ( .A1(\mreg/_02571_ ), .A2(\mreg/_04101_ ), .A3(\mreg/_02566_ ), .ZN(\mreg/_02928_ ) );
NAND3_X1 \mreg/_08840_ ( .A1(\mreg/_02696_ ), .A2(\mreg/_04069_ ), .A3(\mreg/_02633_ ), .ZN(\mreg/_02929_ ) );
NAND3_X1 \mreg/_08841_ ( .A1(\mreg/_02699_ ), .A2(\mreg/_04133_ ), .A3(\mreg/_02691_ ), .ZN(\mreg/_02930_ ) );
AND4_X1 \mreg/_08842_ ( .A1(\mreg/_02927_ ), .A2(\mreg/_02928_ ), .A3(\mreg/_02929_ ), .A4(\mreg/_02930_ ), .ZN(\mreg/_02931_ ) );
AND4_X1 \mreg/_08843_ ( .A1(\mreg/_02917_ ), .A2(\mreg/_02921_ ), .A3(\mreg/_02926_ ), .A4(\mreg/_02931_ ), .ZN(\mreg/_02932_ ) );
NAND4_X1 \mreg/_08844_ ( .A1(\mreg/_02586_ ), .A2(\mreg/_04229_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02579_ ), .ZN(\mreg/_02933_ ) );
OAI21_X1 \mreg/_08845_ ( .A(\mreg/_02933_ ), .B1(\mreg/_02493_ ), .B2(\mreg/_01575_ ), .ZN(\mreg/_02934_ ) );
AOI221_X4 \mreg/_08846_ ( .A(\mreg/_02934_ ), .B1(\mreg/_04197_ ), .B2(\mreg/_02496_ ), .C1(\mreg/_04165_ ), .C2(\mreg/_02501_ ), .ZN(\mreg/_02935_ ) );
NAND3_X1 \mreg/_08847_ ( .A1(\mreg/_02506_ ), .A2(\mreg/_04389_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02936_ ) );
NAND3_X1 \mreg/_08848_ ( .A1(\mreg/_02508_ ), .A2(\mreg/_04421_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02937_ ) );
NAND3_X1 \mreg/_08849_ ( .A1(\mreg/_02503_ ), .A2(\mreg/_04357_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02938_ ) );
NAND3_X1 \mreg/_08850_ ( .A1(\mreg/_02511_ ), .A2(\mreg/_04325_ ), .A3(\mreg/_02513_ ), .ZN(\mreg/_02939_ ) );
AND4_X1 \mreg/_08851_ ( .A1(\mreg/_02936_ ), .A2(\mreg/_02937_ ), .A3(\mreg/_02938_ ), .A4(\mreg/_02939_ ), .ZN(\mreg/_02940_ ) );
NAND4_X1 \mreg/_08852_ ( .A1(\mreg/_02915_ ), .A2(\mreg/_02932_ ), .A3(\mreg/_02935_ ), .A4(\mreg/_02940_ ), .ZN(\mreg/_03909_ ) );
NAND3_X1 \mreg/_08853_ ( .A1(\mreg/_02672_ ), .A2(\mreg/_04359_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02941_ ) );
NAND4_X1 \mreg/_08854_ ( .A1(\mreg/_02535_ ), .A2(\mreg/_04199_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02609_ ), .ZN(\mreg/_02942_ ) );
OAI21_X1 \mreg/_08855_ ( .A(\mreg/_02942_ ), .B1(\mreg/_02493_ ), .B2(\mreg/_01614_ ), .ZN(\mreg/_02943_ ) );
AOI221_X4 \mreg/_08856_ ( .A(\mreg/_02943_ ), .B1(\mreg/_04167_ ), .B2(\mreg/_02496_ ), .C1(\mreg/_04135_ ), .C2(\mreg/_02501_ ), .ZN(\mreg/_02944_ ) );
NAND3_X1 \mreg/_08857_ ( .A1(\mreg/_02674_ ), .A2(\mreg/_04391_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02945_ ) );
AND3_X1 \mreg/_08858_ ( .A1(\mreg/_02619_ ), .A2(\mreg/_04295_ ), .A3(\mreg/_02467_ ), .ZN(\mreg/_02946_ ) );
AND2_X1 \mreg/_08859_ ( .A1(\mreg/_02462_ ), .A2(\mreg/_03872_ ), .ZN(\mreg/_02947_ ) );
AOI21_X1 \mreg/_08860_ ( .A(\mreg/_02946_ ), .B1(\mreg/_04327_ ), .B2(\mreg/_02947_ ), .ZN(\mreg/_02948_ ) );
AND4_X1 \mreg/_08861_ ( .A1(\mreg/_02941_ ), .A2(\mreg/_02944_ ), .A3(\mreg/_02945_ ), .A4(\mreg/_02948_ ), .ZN(\mreg/_02949_ ) );
NAND3_X1 \mreg/_08862_ ( .A1(\mreg/_02531_ ), .A2(\mreg/_04551_ ), .A3(\mreg/_02533_ ), .ZN(\mreg/_02950_ ) );
NAND3_X1 \mreg/_08863_ ( .A1(\mreg/_02516_ ), .A2(\mreg/_04647_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02951_ ) );
NAND3_X1 \mreg/_08864_ ( .A1(\mreg/_02546_ ), .A2(\mreg/_04583_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02952_ ) );
NAND3_X1 \mreg/_08865_ ( .A1(\mreg/_02524_ ), .A2(\mreg/_01601_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02953_ ) );
AND4_X1 \mreg/_08866_ ( .A1(\mreg/_02950_ ), .A2(\mreg/_02951_ ), .A3(\mreg/_02952_ ), .A4(\mreg/_02953_ ), .ZN(\mreg/_02954_ ) );
NAND4_X1 \mreg/_08867_ ( .A1(\mreg/_02586_ ), .A2(\mreg/_02644_ ), .A3(\mreg/_04487_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_02955_ ) );
OAI21_X1 \mreg/_08868_ ( .A(\mreg/_02955_ ), .B1(\mreg/_02539_ ), .B2(\mreg/_01605_ ), .ZN(\mreg/_02956_ ) );
AOI221_X4 \mreg/_08869_ ( .A(\mreg/_02956_ ), .B1(\mreg/_04455_ ), .B2(\mreg/_02542_ ), .C1(\mreg/_04423_ ), .C2(\mreg/_02544_ ), .ZN(\mreg/_02957_ ) );
AND3_X1 \mreg/_08870_ ( .A1(\mreg/_02409_ ), .A2(\mreg/_04615_ ), .A3(\mreg/_02415_ ), .ZN(\mreg/_02958_ ) );
AOI221_X4 \mreg/_08871_ ( .A(\mreg/_02958_ ), .B1(\mreg/_02416_ ), .B2(\mreg/_04711_ ), .C1(\mreg/_04263_ ), .C2(\mreg/_02421_ ), .ZN(\mreg/_02959_ ) );
NAND3_X1 \mreg/_08872_ ( .A1(\mreg/_02463_ ), .A2(\mreg/_04775_ ), .A3(\mreg/_02460_ ), .ZN(\mreg/_02960_ ) );
NAND3_X1 \mreg/_08873_ ( .A1(\mreg/_02454_ ), .A2(\mreg/_04807_ ), .A3(\mreg/_02486_ ), .ZN(\mreg/_02961_ ) );
NAND3_X1 \mreg/_08874_ ( .A1(\mreg/_02632_ ), .A2(\mreg/_04839_ ), .A3(\mreg/_02572_ ), .ZN(\mreg/_02962_ ) );
NAND3_X1 \mreg/_08875_ ( .A1(\mreg/_02684_ ), .A2(\mreg/_02568_ ), .A3(\mreg/_04743_ ), .ZN(\mreg/_02963_ ) );
AND4_X1 \mreg/_08876_ ( .A1(\mreg/_02960_ ), .A2(\mreg/_02961_ ), .A3(\mreg/_02962_ ), .A4(\mreg/_02963_ ), .ZN(\mreg/_02964_ ) );
NAND3_X1 \mreg/_08877_ ( .A1(\mreg/_02471_ ), .A2(\mreg/_04903_ ), .A3(\mreg/_02464_ ), .ZN(\mreg/_02965_ ) );
NAND3_X1 \mreg/_08878_ ( .A1(\mreg/_02476_ ), .A2(\mreg/_03943_ ), .A3(\mreg/_02688_ ), .ZN(\mreg/_02966_ ) );
NAND3_X1 \mreg/_08879_ ( .A1(\mreg/_02684_ ), .A2(\mreg/_02481_ ), .A3(\mreg/_04871_ ), .ZN(\mreg/_02967_ ) );
NAND3_X1 \mreg/_08880_ ( .A1(\mreg/_02485_ ), .A2(\mreg/_03975_ ), .A3(\mreg/_02691_ ), .ZN(\mreg/_02968_ ) );
AND4_X1 \mreg/_08881_ ( .A1(\mreg/_02965_ ), .A2(\mreg/_02966_ ), .A3(\mreg/_02967_ ), .A4(\mreg/_02968_ ), .ZN(\mreg/_02969_ ) );
NAND3_X1 \mreg/_08882_ ( .A1(\mreg/_02479_ ), .A2(\mreg/_04007_ ), .A3(\mreg/_02664_ ), .ZN(\mreg/_02970_ ) );
NAND3_X1 \mreg/_08883_ ( .A1(\mreg/_02431_ ), .A2(\mreg/_04071_ ), .A3(\mreg/_02633_ ), .ZN(\mreg/_02971_ ) );
NAND3_X1 \mreg/_08884_ ( .A1(\mreg/_02440_ ), .A2(\mreg/_04039_ ), .A3(\mreg/_02697_ ), .ZN(\mreg/_02972_ ) );
NAND3_X1 \mreg/_08885_ ( .A1(\mreg/_02699_ ), .A2(\mreg/_04103_ ), .A3(\mreg/_02700_ ), .ZN(\mreg/_02973_ ) );
AND4_X1 \mreg/_08886_ ( .A1(\mreg/_02970_ ), .A2(\mreg/_02971_ ), .A3(\mreg/_02972_ ), .A4(\mreg/_02973_ ), .ZN(\mreg/_02974_ ) );
AND4_X1 \mreg/_08887_ ( .A1(\mreg/_02959_ ), .A2(\mreg/_02964_ ), .A3(\mreg/_02969_ ), .A4(\mreg/_02974_ ), .ZN(\mreg/_02975_ ) );
NAND4_X1 \mreg/_08888_ ( .A1(\mreg/_02949_ ), .A2(\mreg/_02954_ ), .A3(\mreg/_02957_ ), .A4(\mreg/_02975_ ), .ZN(\mreg/_03879_ ) );
NAND3_X1 \mreg/_08889_ ( .A1(\mreg/_02672_ ), .A2(\mreg/_04360_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02976_ ) );
NAND4_X1 \mreg/_08890_ ( .A1(\mreg/_02535_ ), .A2(\mreg/_04200_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02609_ ), .ZN(\mreg/_02977_ ) );
OAI21_X1 \mreg/_08891_ ( .A(\mreg/_02977_ ), .B1(\mreg/_02493_ ), .B2(\mreg/_01669_ ), .ZN(\mreg/_02978_ ) );
AOI221_X4 \mreg/_08892_ ( .A(\mreg/_02978_ ), .B1(\mreg/_04168_ ), .B2(\mreg/_02496_ ), .C1(\mreg/_04136_ ), .C2(\mreg/_02501_ ), .ZN(\mreg/_02979_ ) );
NAND3_X1 \mreg/_08893_ ( .A1(\mreg/_02674_ ), .A2(\mreg/_04392_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02980_ ) );
AND3_X1 \mreg/_08894_ ( .A1(\mreg/_02619_ ), .A2(\mreg/_04296_ ), .A3(\mreg/_02467_ ), .ZN(\mreg/_02981_ ) );
AOI21_X1 \mreg/_08895_ ( .A(\mreg/_02981_ ), .B1(\mreg/_04328_ ), .B2(\mreg/_02947_ ), .ZN(\mreg/_02982_ ) );
AND4_X1 \mreg/_08896_ ( .A1(\mreg/_02976_ ), .A2(\mreg/_02979_ ), .A3(\mreg/_02980_ ), .A4(\mreg/_02982_ ), .ZN(\mreg/_02983_ ) );
AND3_X1 \mreg/_08897_ ( .A1(\mreg/_02597_ ), .A2(\mreg/_04584_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02984_ ) );
AND3_X1 \mreg/_08898_ ( .A1(\mreg/_02599_ ), .A2(\mreg/_04552_ ), .A3(\mreg/_02446_ ), .ZN(\mreg/_02985_ ) );
OR2_X1 \mreg/_08899_ ( .A1(\mreg/_02984_ ), .A2(\mreg/_02985_ ), .ZN(\mreg/_02986_ ) );
AOI221_X4 \mreg/_08900_ ( .A(\mreg/_02986_ ), .B1(\mreg/_01664_ ), .B2(\mreg/_02550_ ), .C1(\mreg/_04648_ ), .C2(\mreg/_02603_ ), .ZN(\mreg/_02987_ ) );
AND3_X1 \mreg/_08901_ ( .A1(\mreg/_02639_ ), .A2(\mreg/_04456_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_02988_ ) );
AND3_X1 \mreg/_08902_ ( .A1(\mreg/_02511_ ), .A2(\mreg/_04424_ ), .A3(\mreg/_02645_ ), .ZN(\mreg/_02989_ ) );
AND4_X1 \mreg/_08903_ ( .A1(\mreg/_04488_ ), .A2(\mreg/_02586_ ), .A3(\mreg/_02851_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_02990_ ) );
AND4_X1 \mreg/_08904_ ( .A1(\mreg/_04520_ ), .A2(\mreg/_02851_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02589_ ), .ZN(\mreg/_02991_ ) );
NOR4_X1 \mreg/_08905_ ( .A1(\mreg/_02988_ ), .A2(\mreg/_02989_ ), .A3(\mreg/_02990_ ), .A4(\mreg/_02991_ ), .ZN(\mreg/_02992_ ) );
AND3_X1 \mreg/_08906_ ( .A1(\mreg/_02855_ ), .A2(\mreg/_04712_ ), .A3(\mreg/_02415_ ), .ZN(\mreg/_02993_ ) );
AOI221_X4 \mreg/_08907_ ( .A(\mreg/_02993_ ), .B1(\mreg/_02627_ ), .B2(\mreg/_04616_ ), .C1(\mreg/_04264_ ), .C2(\mreg/_02421_ ), .ZN(\mreg/_02994_ ) );
NAND3_X1 \mreg/_08908_ ( .A1(\mreg/_02463_ ), .A2(\mreg/_04776_ ), .A3(\mreg/_02460_ ), .ZN(\mreg/_02995_ ) );
NAND3_X1 \mreg/_08909_ ( .A1(\mreg/_02454_ ), .A2(\mreg/_04808_ ), .A3(\mreg/_02486_ ), .ZN(\mreg/_02996_ ) );
NAND3_X1 \mreg/_08910_ ( .A1(\mreg/_02632_ ), .A2(\mreg/_04840_ ), .A3(\mreg/_02572_ ), .ZN(\mreg/_02997_ ) );
NAND3_X1 \mreg/_08911_ ( .A1(\mreg/_02684_ ), .A2(\mreg/_02568_ ), .A3(\mreg/_04744_ ), .ZN(\mreg/_02998_ ) );
AND4_X1 \mreg/_08912_ ( .A1(\mreg/_02995_ ), .A2(\mreg/_02996_ ), .A3(\mreg/_02997_ ), .A4(\mreg/_02998_ ), .ZN(\mreg/_02999_ ) );
NAND3_X1 \mreg/_08913_ ( .A1(\mreg/_02471_ ), .A2(\mreg/_04904_ ), .A3(\mreg/_02464_ ), .ZN(\mreg/_03000_ ) );
NAND3_X1 \mreg/_08914_ ( .A1(\mreg/_02476_ ), .A2(\mreg/_03944_ ), .A3(\mreg/_02688_ ), .ZN(\mreg/_03001_ ) );
NAND3_X1 \mreg/_08915_ ( .A1(\mreg/_02684_ ), .A2(\mreg/_02481_ ), .A3(\mreg/_04872_ ), .ZN(\mreg/_03002_ ) );
NAND3_X1 \mreg/_08916_ ( .A1(\mreg/_02484_ ), .A2(\mreg/_03976_ ), .A3(\mreg/_02691_ ), .ZN(\mreg/_03003_ ) );
AND4_X1 \mreg/_08917_ ( .A1(\mreg/_03000_ ), .A2(\mreg/_03001_ ), .A3(\mreg/_03002_ ), .A4(\mreg/_03003_ ), .ZN(\mreg/_03004_ ) );
NAND3_X1 \mreg/_08918_ ( .A1(\mreg/_02479_ ), .A2(\mreg/_04008_ ), .A3(\mreg/_02664_ ), .ZN(\mreg/_03005_ ) );
NAND3_X1 \mreg/_08919_ ( .A1(\mreg/_02431_ ), .A2(\mreg/_04072_ ), .A3(\mreg/_02633_ ), .ZN(\mreg/_03006_ ) );
NAND3_X1 \mreg/_08920_ ( .A1(\mreg/_02440_ ), .A2(\mreg/_04040_ ), .A3(\mreg/_02697_ ), .ZN(\mreg/_03007_ ) );
NAND3_X1 \mreg/_08921_ ( .A1(\mreg/_02425_ ), .A2(\mreg/_04104_ ), .A3(\mreg/_02700_ ), .ZN(\mreg/_03008_ ) );
AND4_X1 \mreg/_08922_ ( .A1(\mreg/_03005_ ), .A2(\mreg/_03006_ ), .A3(\mreg/_03007_ ), .A4(\mreg/_03008_ ), .ZN(\mreg/_03009_ ) );
AND4_X2 \mreg/_08923_ ( .A1(\mreg/_02994_ ), .A2(\mreg/_02999_ ), .A3(\mreg/_03004_ ), .A4(\mreg/_03009_ ), .ZN(\mreg/_03010_ ) );
NAND4_X1 \mreg/_08924_ ( .A1(\mreg/_02983_ ), .A2(\mreg/_02987_ ), .A3(\mreg/_02992_ ), .A4(\mreg/_03010_ ), .ZN(\mreg/_03880_ ) );
NAND3_X1 \mreg/_08925_ ( .A1(\mreg/_02597_ ), .A2(\mreg/_04585_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03011_ ) );
NAND3_X1 \mreg/_08926_ ( .A1(\mreg/_02599_ ), .A2(\mreg/_04553_ ), .A3(\mreg/_02446_ ), .ZN(\mreg/_03012_ ) );
NAND2_X1 \mreg/_08927_ ( .A1(\mreg/_03011_ ), .A2(\mreg/_03012_ ), .ZN(\mreg/_03013_ ) );
AOI221_X4 \mreg/_08928_ ( .A(\mreg/_03013_ ), .B1(\mreg/_01684_ ), .B2(\mreg/_02549_ ), .C1(\mreg/_04649_ ), .C2(\mreg/_02603_ ), .ZN(\mreg/_03014_ ) );
BUF_X4 \mreg/_08929_ ( .A(\mreg/_02451_ ), .Z(\mreg/_03015_ ) );
NAND4_X1 \mreg/_08930_ ( .A1(\mreg/_03015_ ), .A2(\mreg/_02879_ ), .A3(\mreg/_04489_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03016_ ) );
OAI21_X1 \mreg/_08931_ ( .A(\mreg/_03016_ ), .B1(\mreg/_02660_ ), .B2(\mreg/_01679_ ), .ZN(\mreg/_03017_ ) );
AOI221_X4 \mreg/_08932_ ( .A(\mreg/_03017_ ), .B1(\mreg/_04457_ ), .B2(\mreg/_02759_ ), .C1(\mreg/_04425_ ), .C2(\mreg/_02760_ ), .ZN(\mreg/_03018_ ) );
NAND4_X1 \mreg/_08933_ ( .A1(\mreg/_02608_ ), .A2(\mreg/_04201_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02499_ ), .ZN(\mreg/_03019_ ) );
OAI21_X1 \mreg/_08934_ ( .A(\mreg/_03019_ ), .B1(\mreg/_02611_ ), .B2(\mreg/_01688_ ), .ZN(\mreg/_03020_ ) );
AOI221_X4 \mreg/_08935_ ( .A(\mreg/_03020_ ), .B1(\mreg/_04169_ ), .B2(\mreg/_02613_ ), .C1(\mreg/_04137_ ), .C2(\mreg/_02614_ ), .ZN(\mreg/_03021_ ) );
NAND3_X1 \mreg/_08936_ ( .A1(\mreg/_02715_ ), .A2(\mreg/_04361_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03022_ ) );
NAND3_X1 \mreg/_08937_ ( .A1(\mreg/_02565_ ), .A2(\mreg/_04393_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03023_ ) );
NAND3_X1 \mreg/_08938_ ( .A1(\mreg/_02767_ ), .A2(\mreg/_04329_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03024_ ) );
NAND3_X1 \mreg/_08939_ ( .A1(\mreg/_02520_ ), .A2(\mreg/_04297_ ), .A3(\mreg/_02467_ ), .ZN(\mreg/_03025_ ) );
AND4_X1 \mreg/_08940_ ( .A1(\mreg/_03022_ ), .A2(\mreg/_03023_ ), .A3(\mreg/_03024_ ), .A4(\mreg/_03025_ ), .ZN(\mreg/_03026_ ) );
AND4_X2 \mreg/_08941_ ( .A1(\mreg/_03014_ ), .A2(\mreg/_03018_ ), .A3(\mreg/_03021_ ), .A4(\mreg/_03026_ ), .ZN(\mreg/_03027_ ) );
NAND3_X1 \mreg/_08942_ ( .A1(\mreg/_02583_ ), .A2(\mreg/_04265_ ), .A3(\mreg/_02624_ ), .ZN(\mreg/_03028_ ) );
AND3_X1 \mreg/_08943_ ( .A1(\mreg/_02565_ ), .A2(\mreg/_04841_ ), .A3(\mreg/_02563_ ), .ZN(\mreg/_03029_ ) );
AOI21_X1 \mreg/_08944_ ( .A(\mreg/_03029_ ), .B1(\mreg/_04809_ ), .B2(\mreg/_02636_ ), .ZN(\mreg/_03030_ ) );
AOI22_X1 \mreg/_08945_ ( .A1(\mreg/_04617_ ), .A2(\mreg/_02724_ ), .B1(\mreg/_02723_ ), .B2(\mreg/_04713_ ), .ZN(\mreg/_03031_ ) );
AOI22_X1 \mreg/_08946_ ( .A1(\mreg/_02815_ ), .A2(\mreg/_04777_ ), .B1(\mreg/_04745_ ), .B2(\mreg/_02817_ ), .ZN(\mreg/_03032_ ) );
AND4_X1 \mreg/_08947_ ( .A1(\mreg/_03028_ ), .A2(\mreg/_03030_ ), .A3(\mreg/_03031_ ), .A4(\mreg/_03032_ ), .ZN(\mreg/_03033_ ) );
NAND3_X1 \mreg/_08948_ ( .A1(\mreg/_02639_ ), .A2(\mreg/_04905_ ), .A3(\mreg/_02624_ ), .ZN(\mreg/_03034_ ) );
NAND3_X1 \mreg/_08949_ ( .A1(\mreg/_02641_ ), .A2(\mreg/_03945_ ), .A3(\mreg/_02642_ ), .ZN(\mreg/_03035_ ) );
NAND3_X1 \mreg/_08950_ ( .A1(\mreg/_02630_ ), .A2(\mreg/_02645_ ), .A3(\mreg/_04873_ ), .ZN(\mreg/_03036_ ) );
NAND3_X1 \mreg/_08951_ ( .A1(\mreg/_02647_ ), .A2(\mreg/_03977_ ), .A3(\mreg/_02648_ ), .ZN(\mreg/_03037_ ) );
AND4_X1 \mreg/_08952_ ( .A1(\mreg/_03034_ ), .A2(\mreg/_03035_ ), .A3(\mreg/_03036_ ), .A4(\mreg/_03037_ ), .ZN(\mreg/_03038_ ) );
NAND3_X1 \mreg/_08953_ ( .A1(\mreg/_02630_ ), .A2(\mreg/_04009_ ), .A3(\mreg/_02742_ ), .ZN(\mreg/_03039_ ) );
NAND3_X1 \mreg/_08954_ ( .A1(\mreg/_02785_ ), .A2(\mreg/_04073_ ), .A3(\mreg/_02652_ ), .ZN(\mreg/_03040_ ) );
NAND3_X1 \mreg/_08955_ ( .A1(\mreg/_02744_ ), .A2(\mreg/_04041_ ), .A3(\mreg/_02654_ ), .ZN(\mreg/_03041_ ) );
NAND3_X1 \mreg/_08956_ ( .A1(\mreg/_02787_ ), .A2(\mreg/_04105_ ), .A3(\mreg/_02648_ ), .ZN(\mreg/_03042_ ) );
AND4_X1 \mreg/_08957_ ( .A1(\mreg/_03039_ ), .A2(\mreg/_03040_ ), .A3(\mreg/_03041_ ), .A4(\mreg/_03042_ ), .ZN(\mreg/_03043_ ) );
NAND4_X1 \mreg/_08958_ ( .A1(\mreg/_03027_ ), .A2(\mreg/_03033_ ), .A3(\mreg/_03038_ ), .A4(\mreg/_03043_ ), .ZN(\mreg/_03881_ ) );
NAND3_X1 \mreg/_08959_ ( .A1(\mreg/_02597_ ), .A2(\mreg/_04586_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03044_ ) );
NAND3_X1 \mreg/_08960_ ( .A1(\mreg/_02599_ ), .A2(\mreg/_04554_ ), .A3(\mreg/_02446_ ), .ZN(\mreg/_03045_ ) );
NAND2_X1 \mreg/_08961_ ( .A1(\mreg/_03044_ ), .A2(\mreg/_03045_ ), .ZN(\mreg/_03046_ ) );
AOI221_X4 \mreg/_08962_ ( .A(\mreg/_03046_ ), .B1(\mreg/_01716_ ), .B2(\mreg/_02549_ ), .C1(\mreg/_04650_ ), .C2(\mreg/_02603_ ), .ZN(\mreg/_03047_ ) );
NAND4_X1 \mreg/_08963_ ( .A1(\mreg/_03015_ ), .A2(\mreg/_02879_ ), .A3(\mreg/_04490_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03048_ ) );
OAI21_X1 \mreg/_08964_ ( .A(\mreg/_03048_ ), .B1(\mreg/_02660_ ), .B2(\mreg/_01721_ ), .ZN(\mreg/_03049_ ) );
AOI221_X4 \mreg/_08965_ ( .A(\mreg/_03049_ ), .B1(\mreg/_04458_ ), .B2(\mreg/_02759_ ), .C1(\mreg/_04426_ ), .C2(\mreg/_02760_ ), .ZN(\mreg/_03050_ ) );
NAND4_X1 \mreg/_08966_ ( .A1(\mreg/_02608_ ), .A2(\mreg/_04202_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02499_ ), .ZN(\mreg/_03051_ ) );
OAI21_X1 \mreg/_08967_ ( .A(\mreg/_03051_ ), .B1(\mreg/_02611_ ), .B2(\mreg/_01729_ ), .ZN(\mreg/_03052_ ) );
AOI221_X4 \mreg/_08968_ ( .A(\mreg/_03052_ ), .B1(\mreg/_04170_ ), .B2(\mreg/_02613_ ), .C1(\mreg/_04138_ ), .C2(\mreg/_02614_ ), .ZN(\mreg/_03053_ ) );
NAND3_X1 \mreg/_08969_ ( .A1(\mreg/_02715_ ), .A2(\mreg/_04362_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03054_ ) );
NAND3_X1 \mreg/_08970_ ( .A1(\mreg/_02565_ ), .A2(\mreg/_04394_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03055_ ) );
NAND3_X1 \mreg/_08971_ ( .A1(\mreg/_02767_ ), .A2(\mreg/_04330_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03056_ ) );
NAND3_X1 \mreg/_08972_ ( .A1(\mreg/_02520_ ), .A2(\mreg/_04298_ ), .A3(\mreg/_02467_ ), .ZN(\mreg/_03057_ ) );
AND4_X1 \mreg/_08973_ ( .A1(\mreg/_03054_ ), .A2(\mreg/_03055_ ), .A3(\mreg/_03056_ ), .A4(\mreg/_03057_ ), .ZN(\mreg/_03058_ ) );
AND4_X2 \mreg/_08974_ ( .A1(\mreg/_03047_ ), .A2(\mreg/_03050_ ), .A3(\mreg/_03053_ ), .A4(\mreg/_03058_ ), .ZN(\mreg/_03059_ ) );
NAND3_X1 \mreg/_08975_ ( .A1(\mreg/_02583_ ), .A2(\mreg/_04266_ ), .A3(\mreg/_02624_ ), .ZN(\mreg/_03060_ ) );
AND3_X1 \mreg/_08976_ ( .A1(\mreg/_02565_ ), .A2(\mreg/_04842_ ), .A3(\mreg/_02563_ ), .ZN(\mreg/_03061_ ) );
AOI21_X1 \mreg/_08977_ ( .A(\mreg/_03061_ ), .B1(\mreg/_04810_ ), .B2(\mreg/_02636_ ), .ZN(\mreg/_03062_ ) );
AOI22_X1 \mreg/_08978_ ( .A1(\mreg/_04618_ ), .A2(\mreg/_02724_ ), .B1(\mreg/_02723_ ), .B2(\mreg/_04714_ ), .ZN(\mreg/_03063_ ) );
AOI22_X1 \mreg/_08979_ ( .A1(\mreg/_02815_ ), .A2(\mreg/_04778_ ), .B1(\mreg/_04746_ ), .B2(\mreg/_02817_ ), .ZN(\mreg/_03064_ ) );
AND4_X1 \mreg/_08980_ ( .A1(\mreg/_03060_ ), .A2(\mreg/_03062_ ), .A3(\mreg/_03063_ ), .A4(\mreg/_03064_ ), .ZN(\mreg/_03065_ ) );
NAND3_X1 \mreg/_08981_ ( .A1(\mreg/_02639_ ), .A2(\mreg/_04906_ ), .A3(\mreg/_02820_ ), .ZN(\mreg/_03066_ ) );
NAND3_X1 \mreg/_08982_ ( .A1(\mreg/_02641_ ), .A2(\mreg/_03946_ ), .A3(\mreg/_02642_ ), .ZN(\mreg/_03067_ ) );
NAND3_X1 \mreg/_08983_ ( .A1(\mreg/_02630_ ), .A2(\mreg/_02645_ ), .A3(\mreg/_04874_ ), .ZN(\mreg/_03068_ ) );
NAND3_X1 \mreg/_08984_ ( .A1(\mreg/_02647_ ), .A2(\mreg/_03978_ ), .A3(\mreg/_02648_ ), .ZN(\mreg/_03069_ ) );
AND4_X1 \mreg/_08985_ ( .A1(\mreg/_03066_ ), .A2(\mreg/_03067_ ), .A3(\mreg/_03068_ ), .A4(\mreg/_03069_ ), .ZN(\mreg/_03070_ ) );
NAND3_X1 \mreg/_08986_ ( .A1(\mreg/_02630_ ), .A2(\mreg/_04010_ ), .A3(\mreg/_02742_ ), .ZN(\mreg/_03071_ ) );
NAND3_X1 \mreg/_08987_ ( .A1(\mreg/_02785_ ), .A2(\mreg/_04074_ ), .A3(\mreg/_02652_ ), .ZN(\mreg/_03072_ ) );
NAND3_X1 \mreg/_08988_ ( .A1(\mreg/_02744_ ), .A2(\mreg/_04042_ ), .A3(\mreg/_02654_ ), .ZN(\mreg/_03073_ ) );
NAND3_X1 \mreg/_08989_ ( .A1(\mreg/_02787_ ), .A2(\mreg/_04106_ ), .A3(\mreg/_02648_ ), .ZN(\mreg/_03074_ ) );
AND4_X1 \mreg/_08990_ ( .A1(\mreg/_03071_ ), .A2(\mreg/_03072_ ), .A3(\mreg/_03073_ ), .A4(\mreg/_03074_ ), .ZN(\mreg/_03075_ ) );
NAND4_X1 \mreg/_08991_ ( .A1(\mreg/_03059_ ), .A2(\mreg/_03065_ ), .A3(\mreg/_03070_ ), .A4(\mreg/_03075_ ), .ZN(\mreg/_03882_ ) );
NAND3_X1 \mreg/_08992_ ( .A1(\mreg/_02855_ ), .A2(\mreg/_04715_ ), .A3(\mreg/_02411_ ), .ZN(\mreg/_03076_ ) );
NAND3_X1 \mreg/_08993_ ( .A1(\mreg/_02443_ ), .A2(\mreg/_02452_ ), .A3(\mreg/_04747_ ), .ZN(\mreg/_03077_ ) );
NAND2_X1 \mreg/_08994_ ( .A1(\mreg/_03076_ ), .A2(\mreg/_03077_ ), .ZN(\mreg/_03078_ ) );
AOI221_X4 \mreg/_08995_ ( .A(\mreg/_03078_ ), .B1(\mreg/_04779_ ), .B2(\mreg/_02814_ ), .C1(\mreg/_04811_ ), .C2(\mreg/_02635_ ), .ZN(\mreg/_03079_ ) );
NAND4_X1 \mreg/_08996_ ( .A1(\mreg/_03015_ ), .A2(\mreg/_02879_ ), .A3(\mreg/_04491_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03080_ ) );
OAI21_X1 \mreg/_08997_ ( .A(\mreg/_03080_ ), .B1(\mreg/_02660_ ), .B2(\mreg/_01755_ ), .ZN(\mreg/_03081_ ) );
AOI221_X4 \mreg/_08998_ ( .A(\mreg/_03081_ ), .B1(\mreg/_01752_ ), .B2(\mreg/_02549_ ), .C1(\mreg/_04651_ ), .C2(\mreg/_02603_ ), .ZN(\mreg/_03082_ ) );
NAND3_X1 \mreg/_08999_ ( .A1(\mreg/_02597_ ), .A2(\mreg/_04043_ ), .A3(\mreg/_02553_ ), .ZN(\mreg/_03083_ ) );
NAND3_X1 \mreg/_09000_ ( .A1(\mreg/_02424_ ), .A2(\mreg/_04107_ ), .A3(\mreg/_02553_ ), .ZN(\mreg/_03084_ ) );
NAND2_X1 \mreg/_09001_ ( .A1(\mreg/_03083_ ), .A2(\mreg/_03084_ ), .ZN(\mreg/_03085_ ) );
AOI221_X4 \mreg/_09002_ ( .A(\mreg/_03085_ ), .B1(\mreg/_03947_ ), .B2(\mreg/_02560_ ), .C1(\mreg/_04907_ ), .C2(\mreg/_02734_ ), .ZN(\mreg/_03086_ ) );
NAND3_X1 \mreg/_09003_ ( .A1(\mreg/_02503_ ), .A2(\mreg/_04331_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03087_ ) );
NAND3_X1 \mreg/_09004_ ( .A1(\mreg/_02619_ ), .A2(\mreg/_04299_ ), .A3(\mreg/_02512_ ), .ZN(\mreg/_03088_ ) );
NAND4_X1 \mreg/_09005_ ( .A1(\mreg/_02586_ ), .A2(\mreg/_04203_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02580_ ), .ZN(\mreg/_03089_ ) );
NAND4_X1 \mreg/_09006_ ( .A1(\mreg/_02589_ ), .A2(\mreg/_02580_ ), .A3(\mreg/_04235_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03090_ ) );
AND4_X1 \mreg/_09007_ ( .A1(\mreg/_03087_ ), .A2(\mreg/_03088_ ), .A3(\mreg/_03089_ ), .A4(\mreg/_03090_ ), .ZN(\mreg/_03091_ ) );
AND4_X4 \mreg/_09008_ ( .A1(\mreg/_03079_ ), .A2(\mreg/_03082_ ), .A3(\mreg/_03086_ ), .A4(\mreg/_03091_ ), .ZN(\mreg/_03092_ ) );
NAND3_X1 \mreg/_09009_ ( .A1(\mreg/_02842_ ), .A2(\mreg/_04843_ ), .A3(\mreg/_02779_ ), .ZN(\mreg/_03093_ ) );
NAND3_X1 \mreg/_09010_ ( .A1(\mreg/_02845_ ), .A2(\mreg/_04267_ ), .A3(\mreg/_02779_ ), .ZN(\mreg/_03094_ ) );
NAND3_X1 \mreg/_09011_ ( .A1(\mreg/_02490_ ), .A2(\mreg/_04619_ ), .A3(\mreg/_02779_ ), .ZN(\mreg/_03095_ ) );
NAND3_X1 \mreg/_09012_ ( .A1(\mreg/_02730_ ), .A2(\mreg/_02645_ ), .A3(\mreg/_04875_ ), .ZN(\mreg/_03096_ ) );
NAND4_X1 \mreg/_09013_ ( .A1(\mreg/_03093_ ), .A2(\mreg/_03094_ ), .A3(\mreg/_03095_ ), .A4(\mreg/_03096_ ), .ZN(\mreg/_03097_ ) );
AND3_X1 \mreg/_09014_ ( .A1(\mreg/_02730_ ), .A2(\mreg/_04011_ ), .A3(\mreg/_02742_ ), .ZN(\mreg/_03098_ ) );
AND3_X1 \mreg/_09015_ ( .A1(\mreg/_02485_ ), .A2(\mreg/_03979_ ), .A3(\mreg/_02737_ ), .ZN(\mreg/_03099_ ) );
AND3_X1 \mreg/_09016_ ( .A1(\mreg/_02785_ ), .A2(\mreg/_04075_ ), .A3(\mreg/_02745_ ), .ZN(\mreg/_03100_ ) );
NOR4_X1 \mreg/_09017_ ( .A1(\mreg/_03097_ ), .A2(\mreg/_03098_ ), .A3(\mreg/_03099_ ), .A4(\mreg/_03100_ ), .ZN(\mreg/_03101_ ) );
NAND3_X1 \mreg/_09018_ ( .A1(\mreg/_02696_ ), .A2(\mreg/_04587_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03102_ ) );
NAND3_X1 \mreg/_09019_ ( .A1(\mreg/_02510_ ), .A2(\mreg/_04555_ ), .A3(\mreg/_02447_ ), .ZN(\mreg/_03103_ ) );
NAND2_X1 \mreg/_09020_ ( .A1(\mreg/_03102_ ), .A2(\mreg/_03103_ ), .ZN(\mreg/_03104_ ) );
AOI221_X4 \mreg/_09021_ ( .A(\mreg/_03104_ ), .B1(\mreg/_04459_ ), .B2(\mreg/_02542_ ), .C1(\mreg/_04427_ ), .C2(\mreg/_02544_ ), .ZN(\mreg/_03105_ ) );
NAND3_X1 \mreg/_09022_ ( .A1(\mreg/_02511_ ), .A2(\mreg/_04139_ ), .A3(\mreg/_02581_ ), .ZN(\mreg/_03106_ ) );
NAND3_X1 \mreg/_09023_ ( .A1(\mreg/_02506_ ), .A2(\mreg/_04363_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03107_ ) );
NAND3_X1 \mreg/_09024_ ( .A1(\mreg/_02583_ ), .A2(\mreg/_04171_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03108_ ) );
NAND3_X1 \mreg/_09025_ ( .A1(\mreg/_02508_ ), .A2(\mreg/_04395_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03109_ ) );
AND4_X1 \mreg/_09026_ ( .A1(\mreg/_03106_ ), .A2(\mreg/_03107_ ), .A3(\mreg/_03108_ ), .A4(\mreg/_03109_ ), .ZN(\mreg/_03110_ ) );
NAND4_X1 \mreg/_09027_ ( .A1(\mreg/_03092_ ), .A2(\mreg/_03101_ ), .A3(\mreg/_03105_ ), .A4(\mreg/_03110_ ), .ZN(\mreg/_03883_ ) );
NAND3_X1 \mreg/_09028_ ( .A1(\mreg/_02729_ ), .A2(\mreg/_02466_ ), .A3(\mreg/_04748_ ), .ZN(\mreg/_03111_ ) );
INV_X1 \mreg/_09029_ ( .A(\mreg/_02416_ ), .ZN(\mreg/_03112_ ) );
OAI21_X1 \mreg/_09030_ ( .A(\mreg/_03111_ ), .B1(\mreg/_03112_ ), .B2(\mreg/_01787_ ), .ZN(\mreg/_03113_ ) );
AOI221_X4 \mreg/_09031_ ( .A(\mreg/_03113_ ), .B1(\mreg/_04812_ ), .B2(\mreg/_02635_ ), .C1(\mreg/_04780_ ), .C2(\mreg/_02815_ ), .ZN(\mreg/_03114_ ) );
NAND3_X1 \mreg/_09032_ ( .A1(\mreg/_02425_ ), .A2(\mreg/_04108_ ), .A3(\mreg/_02700_ ), .ZN(\mreg/_03115_ ) );
NAND2_X1 \mreg/_09033_ ( .A1(\mreg/_02440_ ), .A2(\mreg/_02427_ ), .ZN(\mreg/_03116_ ) );
OAI21_X1 \mreg/_09034_ ( .A(\mreg/_03115_ ), .B1(\mreg/_03116_ ), .B2(\mreg/_01792_ ), .ZN(\mreg/_03117_ ) );
AOI221_X4 \mreg/_09035_ ( .A(\mreg/_03117_ ), .B1(\mreg/_03948_ ), .B2(\mreg/_02560_ ), .C1(\mreg/_04908_ ), .C2(\mreg/_02735_ ), .ZN(\mreg/_03118_ ) );
NAND3_X1 \mreg/_09036_ ( .A1(\mreg/_02785_ ), .A2(\mreg/_04652_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03119_ ) );
NAND3_X1 \mreg/_09037_ ( .A1(\mreg/_02787_ ), .A2(\mreg/_01798_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03120_ ) );
NAND4_X1 \mreg/_09038_ ( .A1(\mreg/_02587_ ), .A2(\mreg/_02838_ ), .A3(\mreg/_04492_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03121_ ) );
NAND4_X1 \mreg/_09039_ ( .A1(\mreg/_02645_ ), .A2(\mreg/_04524_ ), .A3(\mreg/_02589_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03122_ ) );
NAND4_X1 \mreg/_09040_ ( .A1(\mreg/_03119_ ), .A2(\mreg/_03120_ ), .A3(\mreg/_03121_ ), .A4(\mreg/_03122_ ), .ZN(\mreg/_03123_ ) );
NAND4_X1 \mreg/_09041_ ( .A1(\mreg/_02587_ ), .A2(\mreg/_04204_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02581_ ), .ZN(\mreg/_03124_ ) );
OAI21_X1 \mreg/_09042_ ( .A(\mreg/_03124_ ), .B1(\mreg/_02493_ ), .B2(\mreg/_01801_ ), .ZN(\mreg/_03125_ ) );
AND3_X1 \mreg/_09043_ ( .A1(\mreg/_02503_ ), .A2(\mreg/_04332_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03126_ ) );
AND3_X1 \mreg/_09044_ ( .A1(\mreg/_02837_ ), .A2(\mreg/_04300_ ), .A3(\mreg/_02512_ ), .ZN(\mreg/_03127_ ) );
NOR4_X1 \mreg/_09045_ ( .A1(\mreg/_03123_ ), .A2(\mreg/_03125_ ), .A3(\mreg/_03126_ ), .A4(\mreg/_03127_ ), .ZN(\mreg/_03128_ ) );
NAND3_X1 \mreg/_09046_ ( .A1(\mreg/_02741_ ), .A2(\mreg/_04012_ ), .A3(\mreg/_02742_ ), .ZN(\mreg/_03129_ ) );
OAI221_X1 \mreg/_09047_ ( .A(\mreg/_03129_ ), .B1(\mreg/_02749_ ), .B2(\mreg/_01806_ ), .C1(\mreg/_01807_ ), .C2(\mreg/_02739_ ), .ZN(\mreg/_03130_ ) );
NAND3_X1 \mreg/_09048_ ( .A1(\mreg/_02472_ ), .A2(\mreg/_04460_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03131_ ) );
NAND3_X1 \mreg/_09049_ ( .A1(\mreg/_02744_ ), .A2(\mreg/_04588_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03132_ ) );
NAND3_X1 \mreg/_09050_ ( .A1(\mreg/_02837_ ), .A2(\mreg/_04556_ ), .A3(\mreg/_02532_ ), .ZN(\mreg/_03133_ ) );
NAND3_X1 \mreg/_09051_ ( .A1(\mreg/_02837_ ), .A2(\mreg/_04428_ ), .A3(\mreg/_02838_ ), .ZN(\mreg/_03134_ ) );
NAND4_X1 \mreg/_09052_ ( .A1(\mreg/_03131_ ), .A2(\mreg/_03132_ ), .A3(\mreg/_03133_ ), .A4(\mreg/_03134_ ), .ZN(\mreg/_03135_ ) );
NAND3_X1 \mreg/_09053_ ( .A1(\mreg/_02455_ ), .A2(\mreg/_04364_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03136_ ) );
NAND3_X1 \mreg/_09054_ ( .A1(\mreg/_02459_ ), .A2(\mreg/_04396_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03137_ ) );
NAND3_X1 \mreg/_09055_ ( .A1(\mreg/_02530_ ), .A2(\mreg/_04140_ ), .A3(\mreg/_02580_ ), .ZN(\mreg/_03138_ ) );
NAND3_X1 \mreg/_09056_ ( .A1(\mreg/_02419_ ), .A2(\mreg/_04172_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03139_ ) );
NAND4_X1 \mreg/_09057_ ( .A1(\mreg/_03136_ ), .A2(\mreg/_03137_ ), .A3(\mreg/_03138_ ), .A4(\mreg/_03139_ ), .ZN(\mreg/_03140_ ) );
NAND3_X1 \mreg/_09058_ ( .A1(\mreg/_02842_ ), .A2(\mreg/_04844_ ), .A3(\mreg/_02747_ ), .ZN(\mreg/_03141_ ) );
NAND3_X1 \mreg/_09059_ ( .A1(\mreg/_02845_ ), .A2(\mreg/_04268_ ), .A3(\mreg/_02623_ ), .ZN(\mreg/_03142_ ) );
NAND3_X1 \mreg/_09060_ ( .A1(\mreg/_02490_ ), .A2(\mreg/_04620_ ), .A3(\mreg/_02623_ ), .ZN(\mreg/_03143_ ) );
NAND3_X1 \mreg/_09061_ ( .A1(\mreg/_02629_ ), .A2(\mreg/_02851_ ), .A3(\mreg/_04876_ ), .ZN(\mreg/_03144_ ) );
NAND4_X1 \mreg/_09062_ ( .A1(\mreg/_03141_ ), .A2(\mreg/_03142_ ), .A3(\mreg/_03143_ ), .A4(\mreg/_03144_ ), .ZN(\mreg/_03145_ ) );
NOR4_X1 \mreg/_09063_ ( .A1(\mreg/_03130_ ), .A2(\mreg/_03135_ ), .A3(\mreg/_03140_ ), .A4(\mreg/_03145_ ), .ZN(\mreg/_03146_ ) );
NAND4_X1 \mreg/_09064_ ( .A1(\mreg/_03114_ ), .A2(\mreg/_03118_ ), .A3(\mreg/_03128_ ), .A4(\mreg/_03146_ ), .ZN(\mreg/_03884_ ) );
NAND3_X1 \mreg/_09065_ ( .A1(\mreg/_02729_ ), .A2(\mreg/_02466_ ), .A3(\mreg/_04749_ ), .ZN(\mreg/_03147_ ) );
OAI21_X1 \mreg/_09066_ ( .A(\mreg/_03147_ ), .B1(\mreg/_03112_ ), .B2(\mreg/_01825_ ), .ZN(\mreg/_03148_ ) );
AOI221_X4 \mreg/_09067_ ( .A(\mreg/_03148_ ), .B1(\mreg/_04813_ ), .B2(\mreg/_02635_ ), .C1(\mreg/_04781_ ), .C2(\mreg/_02815_ ), .ZN(\mreg/_03149_ ) );
AND3_X1 \mreg/_09068_ ( .A1(\mreg/_02462_ ), .A2(\mreg/_04333_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03150_ ) );
AND3_X1 \mreg/_09069_ ( .A1(\mreg/_02510_ ), .A2(\mreg/_04301_ ), .A3(\mreg/_02466_ ), .ZN(\mreg/_03151_ ) );
AND4_X1 \mreg/_09070_ ( .A1(\mreg/_04205_ ), .A2(\mreg/_02585_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02579_ ), .ZN(\mreg/_03152_ ) );
AND4_X1 \mreg/_09071_ ( .A1(\mreg/_04237_ ), .A2(\mreg/_02589_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02579_ ), .ZN(\mreg/_03153_ ) );
OR4_X1 \mreg/_09072_ ( .A1(\mreg/_03150_ ), .A2(\mreg/_03151_ ), .A3(\mreg/_03152_ ), .A4(\mreg/_03153_ ), .ZN(\mreg/_03154_ ) );
AND3_X1 \mreg/_09073_ ( .A1(\mreg/_02785_ ), .A2(\mreg/_04653_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03155_ ) );
AND3_X1 \mreg/_09074_ ( .A1(\mreg/_02787_ ), .A2(\mreg/_01835_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03156_ ) );
NAND4_X1 \mreg/_09075_ ( .A1(\mreg/_02586_ ), .A2(\mreg/_02851_ ), .A3(\mreg/_04493_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03157_ ) );
OAI21_X1 \mreg/_09076_ ( .A(\mreg/_03157_ ), .B1(\mreg/_02539_ ), .B2(\mreg/_01833_ ), .ZN(\mreg/_03158_ ) );
NOR4_X1 \mreg/_09077_ ( .A1(\mreg/_03154_ ), .A2(\mreg/_03155_ ), .A3(\mreg/_03156_ ), .A4(\mreg/_03158_ ), .ZN(\mreg/_03159_ ) );
NAND3_X1 \mreg/_09078_ ( .A1(\mreg/_02425_ ), .A2(\mreg/_04109_ ), .A3(\mreg/_02700_ ), .ZN(\mreg/_03160_ ) );
OAI21_X1 \mreg/_09079_ ( .A(\mreg/_03160_ ), .B1(\mreg/_03116_ ), .B2(\mreg/_01829_ ), .ZN(\mreg/_03161_ ) );
AOI221_X4 \mreg/_09080_ ( .A(\mreg/_03161_ ), .B1(\mreg/_03949_ ), .B2(\mreg/_02560_ ), .C1(\mreg/_04909_ ), .C2(\mreg/_02735_ ), .ZN(\mreg/_03162_ ) );
NAND3_X1 \mreg/_09081_ ( .A1(\mreg/_02741_ ), .A2(\mreg/_04013_ ), .A3(\mreg/_02742_ ), .ZN(\mreg/_03163_ ) );
OAI221_X1 \mreg/_09082_ ( .A(\mreg/_03163_ ), .B1(\mreg/_02749_ ), .B2(\mreg/_01848_ ), .C1(\mreg/_01849_ ), .C2(\mreg/_02739_ ), .ZN(\mreg/_03164_ ) );
NAND3_X1 \mreg/_09083_ ( .A1(\mreg/_02472_ ), .A2(\mreg/_04461_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03165_ ) );
NAND3_X1 \mreg/_09084_ ( .A1(\mreg/_02441_ ), .A2(\mreg/_04589_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03166_ ) );
NAND3_X1 \mreg/_09085_ ( .A1(\mreg/_02837_ ), .A2(\mreg/_04557_ ), .A3(\mreg/_02532_ ), .ZN(\mreg/_03167_ ) );
NAND3_X1 \mreg/_09086_ ( .A1(\mreg/_02530_ ), .A2(\mreg/_04429_ ), .A3(\mreg/_02851_ ), .ZN(\mreg/_03168_ ) );
NAND4_X1 \mreg/_09087_ ( .A1(\mreg/_03165_ ), .A2(\mreg/_03166_ ), .A3(\mreg/_03167_ ), .A4(\mreg/_03168_ ), .ZN(\mreg/_03169_ ) );
NAND3_X1 \mreg/_09088_ ( .A1(\mreg/_02455_ ), .A2(\mreg/_04365_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03170_ ) );
NAND3_X1 \mreg/_09089_ ( .A1(\mreg/_02459_ ), .A2(\mreg/_04397_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03171_ ) );
NAND3_X1 \mreg/_09090_ ( .A1(\mreg/_02530_ ), .A2(\mreg/_04141_ ), .A3(\mreg/_02580_ ), .ZN(\mreg/_03172_ ) );
NAND3_X1 \mreg/_09091_ ( .A1(\mreg/_02419_ ), .A2(\mreg/_04173_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03173_ ) );
NAND4_X1 \mreg/_09092_ ( .A1(\mreg/_03170_ ), .A2(\mreg/_03171_ ), .A3(\mreg/_03172_ ), .A4(\mreg/_03173_ ), .ZN(\mreg/_03174_ ) );
NAND3_X1 \mreg/_09093_ ( .A1(\mreg/_02459_ ), .A2(\mreg/_04845_ ), .A3(\mreg/_02747_ ), .ZN(\mreg/_03175_ ) );
NAND3_X1 \mreg/_09094_ ( .A1(\mreg/_02845_ ), .A2(\mreg/_04269_ ), .A3(\mreg/_02623_ ), .ZN(\mreg/_03176_ ) );
NAND3_X1 \mreg/_09095_ ( .A1(\mreg/_02490_ ), .A2(\mreg/_04621_ ), .A3(\mreg/_02623_ ), .ZN(\mreg/_03177_ ) );
NAND3_X1 \mreg/_09096_ ( .A1(\mreg/_02629_ ), .A2(\mreg/_02851_ ), .A3(\mreg/_04877_ ), .ZN(\mreg/_03178_ ) );
NAND4_X1 \mreg/_09097_ ( .A1(\mreg/_03175_ ), .A2(\mreg/_03176_ ), .A3(\mreg/_03177_ ), .A4(\mreg/_03178_ ), .ZN(\mreg/_03179_ ) );
NOR4_X1 \mreg/_09098_ ( .A1(\mreg/_03164_ ), .A2(\mreg/_03169_ ), .A3(\mreg/_03174_ ), .A4(\mreg/_03179_ ), .ZN(\mreg/_03180_ ) );
NAND4_X1 \mreg/_09099_ ( .A1(\mreg/_03149_ ), .A2(\mreg/_03159_ ), .A3(\mreg/_03162_ ), .A4(\mreg/_03180_ ), .ZN(\mreg/_03885_ ) );
NAND3_X1 \mreg/_09100_ ( .A1(\mreg/_02531_ ), .A2(\mreg/_04558_ ), .A3(\mreg/_02533_ ), .ZN(\mreg/_03181_ ) );
NAND4_X1 \mreg/_09101_ ( .A1(\mreg/_03015_ ), .A2(\mreg/_02879_ ), .A3(\mreg/_04494_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03182_ ) );
OAI21_X1 \mreg/_09102_ ( .A(\mreg/_03182_ ), .B1(\mreg/_02660_ ), .B2(\mreg/_01867_ ), .ZN(\mreg/_03183_ ) );
AOI221_X4 \mreg/_09103_ ( .A(\mreg/_03183_ ), .B1(\mreg/_04462_ ), .B2(\mreg/_02759_ ), .C1(\mreg/_04430_ ), .C2(\mreg/_02760_ ), .ZN(\mreg/_03184_ ) );
NAND3_X1 \mreg/_09104_ ( .A1(\mreg/_02546_ ), .A2(\mreg/_04590_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03185_ ) );
AND3_X1 \mreg/_09105_ ( .A1(\mreg/_02571_ ), .A2(\mreg/_04654_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03186_ ) );
AOI21_X1 \mreg/_09106_ ( .A(\mreg/_03186_ ), .B1(\mreg/_01863_ ), .B2(\mreg/_02550_ ), .ZN(\mreg/_03187_ ) );
AND4_X4 \mreg/_09107_ ( .A1(\mreg/_03181_ ), .A2(\mreg/_03184_ ), .A3(\mreg/_03185_ ), .A4(\mreg/_03187_ ), .ZN(\mreg/_03188_ ) );
NAND3_X1 \mreg/_09108_ ( .A1(\mreg/_02672_ ), .A2(\mreg/_04366_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03189_ ) );
NAND4_X1 \mreg/_09109_ ( .A1(\mreg/_02608_ ), .A2(\mreg/_04206_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02499_ ), .ZN(\mreg/_03190_ ) );
OAI21_X1 \mreg/_09110_ ( .A(\mreg/_03190_ ), .B1(\mreg/_02611_ ), .B2(\mreg/_01875_ ), .ZN(\mreg/_03191_ ) );
AOI221_X4 \mreg/_09111_ ( .A(\mreg/_03191_ ), .B1(\mreg/_04174_ ), .B2(\mreg/_02613_ ), .C1(\mreg/_04142_ ), .C2(\mreg/_02500_ ), .ZN(\mreg/_03192_ ) );
NAND3_X1 \mreg/_09112_ ( .A1(\mreg/_02674_ ), .A2(\mreg/_04398_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03193_ ) );
AND3_X1 \mreg/_09113_ ( .A1(\mreg/_02767_ ), .A2(\mreg/_04334_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03194_ ) );
AOI21_X1 \mreg/_09114_ ( .A(\mreg/_03194_ ), .B1(\mreg/_04302_ ), .B2(\mreg/_02807_ ), .ZN(\mreg/_03195_ ) );
AND4_X1 \mreg/_09115_ ( .A1(\mreg/_03189_ ), .A2(\mreg/_03192_ ), .A3(\mreg/_03193_ ), .A4(\mreg/_03195_ ), .ZN(\mreg/_03196_ ) );
NAND3_X1 \mreg/_09116_ ( .A1(\mreg/_02583_ ), .A2(\mreg/_04270_ ), .A3(\mreg/_02820_ ), .ZN(\mreg/_03197_ ) );
AND3_X1 \mreg/_09117_ ( .A1(\mreg/_02632_ ), .A2(\mreg/_04846_ ), .A3(\mreg/_02566_ ), .ZN(\mreg/_03198_ ) );
AOI21_X1 \mreg/_09118_ ( .A(\mreg/_03198_ ), .B1(\mreg/_04814_ ), .B2(\mreg/_02636_ ), .ZN(\mreg/_03199_ ) );
AOI22_X1 \mreg/_09119_ ( .A1(\mreg/_04622_ ), .A2(\mreg/_02724_ ), .B1(\mreg/_02723_ ), .B2(\mreg/_04718_ ), .ZN(\mreg/_03200_ ) );
AOI22_X1 \mreg/_09120_ ( .A1(\mreg/_02815_ ), .A2(\mreg/_04782_ ), .B1(\mreg/_04750_ ), .B2(\mreg/_02817_ ), .ZN(\mreg/_03201_ ) );
AND4_X1 \mreg/_09121_ ( .A1(\mreg/_03197_ ), .A2(\mreg/_03199_ ), .A3(\mreg/_03200_ ), .A4(\mreg/_03201_ ), .ZN(\mreg/_03202_ ) );
NAND3_X1 \mreg/_09122_ ( .A1(\mreg/_02641_ ), .A2(\mreg/_03950_ ), .A3(\mreg/_02642_ ), .ZN(\mreg/_03203_ ) );
NAND3_X1 \mreg/_09123_ ( .A1(\mreg/_02629_ ), .A2(\mreg/_04014_ ), .A3(\mreg/_02448_ ), .ZN(\mreg/_03204_ ) );
NAND3_X1 \mreg/_09124_ ( .A1(\mreg/_02571_ ), .A2(\mreg/_04078_ ), .A3(\mreg/_02486_ ), .ZN(\mreg/_03205_ ) );
NAND3_X1 \mreg/_09125_ ( .A1(\mreg/_02696_ ), .A2(\mreg/_04046_ ), .A3(\mreg/_02572_ ), .ZN(\mreg/_03206_ ) );
NAND3_X1 \mreg/_09126_ ( .A1(\mreg/_02699_ ), .A2(\mreg/_04110_ ), .A3(\mreg/_02633_ ), .ZN(\mreg/_03207_ ) );
AND4_X1 \mreg/_09127_ ( .A1(\mreg/_03204_ ), .A2(\mreg/_03205_ ), .A3(\mreg/_03206_ ), .A4(\mreg/_03207_ ), .ZN(\mreg/_03208_ ) );
NAND3_X1 \mreg/_09128_ ( .A1(\mreg/_02647_ ), .A2(\mreg/_03982_ ), .A3(\mreg/_02654_ ), .ZN(\mreg/_03209_ ) );
AND3_X1 \mreg/_09129_ ( .A1(\mreg/_02729_ ), .A2(\mreg/_04878_ ), .A3(\mreg/_02644_ ), .ZN(\mreg/_03210_ ) );
AOI21_X1 \mreg/_09130_ ( .A(\mreg/_03210_ ), .B1(\mreg/_02735_ ), .B2(\mreg/_04910_ ), .ZN(\mreg/_03211_ ) );
AND4_X1 \mreg/_09131_ ( .A1(\mreg/_03203_ ), .A2(\mreg/_03208_ ), .A3(\mreg/_03209_ ), .A4(\mreg/_03211_ ), .ZN(\mreg/_03212_ ) );
NAND4_X1 \mreg/_09132_ ( .A1(\mreg/_03188_ ), .A2(\mreg/_03196_ ), .A3(\mreg/_03202_ ), .A4(\mreg/_03212_ ), .ZN(\mreg/_03886_ ) );
NAND4_X1 \mreg/_09133_ ( .A1(\mreg/_02451_ ), .A2(\mreg/_02474_ ), .A3(\mreg/_04495_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03213_ ) );
OAI21_X1 \mreg/_09134_ ( .A(\mreg/_03213_ ), .B1(\mreg/_02538_ ), .B2(\mreg/_01915_ ), .ZN(\mreg/_03214_ ) );
AOI221_X2 \mreg/_09135_ ( .A(\mreg/_03214_ ), .B1(\mreg/_04463_ ), .B2(\mreg/_02541_ ), .C1(\mreg/_04431_ ), .C2(\mreg/_02543_ ), .ZN(\mreg/_03215_ ) );
NAND4_X1 \mreg/_09136_ ( .A1(\mreg/_02451_ ), .A2(\mreg/_04207_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02499_ ), .ZN(\mreg/_03216_ ) );
OAI21_X1 \mreg/_09137_ ( .A(\mreg/_03216_ ), .B1(\mreg/_02492_ ), .B2(\mreg/_01924_ ), .ZN(\mreg/_03217_ ) );
AOI221_X4 \mreg/_09138_ ( .A(\mreg/_03217_ ), .B1(\mreg/_04175_ ), .B2(\mreg/_02495_ ), .C1(\mreg/_04143_ ), .C2(\mreg/_02500_ ), .ZN(\mreg/_03218_ ) );
NAND3_X1 \mreg/_09139_ ( .A1(\mreg/_02597_ ), .A2(\mreg/_04591_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03219_ ) );
NAND3_X1 \mreg/_09140_ ( .A1(\mreg/_02599_ ), .A2(\mreg/_04559_ ), .A3(\mreg/_02446_ ), .ZN(\mreg/_03220_ ) );
NAND2_X1 \mreg/_09141_ ( .A1(\mreg/_03219_ ), .A2(\mreg/_03220_ ), .ZN(\mreg/_03221_ ) );
AOI221_X4 \mreg/_09142_ ( .A(\mreg/_03221_ ), .B1(\mreg/_01920_ ), .B2(\mreg/_02549_ ), .C1(\mreg/_04655_ ), .C2(\mreg/_02602_ ), .ZN(\mreg/_03222_ ) );
NAND3_X1 \mreg/_09143_ ( .A1(\mreg/_02454_ ), .A2(\mreg/_04367_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03223_ ) );
NAND3_X1 \mreg/_09144_ ( .A1(\mreg/_02458_ ), .A2(\mreg/_04399_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03224_ ) );
NAND3_X1 \mreg/_09145_ ( .A1(\mreg/_02462_ ), .A2(\mreg/_04335_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03225_ ) );
NAND3_X1 \mreg/_09146_ ( .A1(\mreg/_02510_ ), .A2(\mreg/_04303_ ), .A3(\mreg/_02466_ ), .ZN(\mreg/_03226_ ) );
AND4_X1 \mreg/_09147_ ( .A1(\mreg/_03223_ ), .A2(\mreg/_03224_ ), .A3(\mreg/_03225_ ), .A4(\mreg/_03226_ ), .ZN(\mreg/_03227_ ) );
NAND4_X1 \mreg/_09148_ ( .A1(\mreg/_03215_ ), .A2(\mreg/_03218_ ), .A3(\mreg/_03222_ ), .A4(\mreg/_03227_ ), .ZN(\mreg/_03228_ ) );
AND3_X1 \mreg/_09149_ ( .A1(\mreg/_02458_ ), .A2(\mreg/_04847_ ), .A3(\mreg/_02427_ ), .ZN(\mreg/_03229_ ) );
AOI21_X1 \mreg/_09150_ ( .A(\mreg/_03229_ ), .B1(\mreg/_04815_ ), .B2(\mreg/_02635_ ), .ZN(\mreg/_03230_ ) );
AOI22_X1 \mreg/_09151_ ( .A1(\mreg/_04623_ ), .A2(\mreg/_02724_ ), .B1(\mreg/_02723_ ), .B2(\mreg/_04719_ ), .ZN(\mreg/_03231_ ) );
NAND3_X1 \mreg/_09152_ ( .A1(\mreg/_02845_ ), .A2(\mreg/_04271_ ), .A3(\mreg/_02737_ ), .ZN(\mreg/_03232_ ) );
AOI22_X1 \mreg/_09153_ ( .A1(\mreg/_02814_ ), .A2(\mreg/_04783_ ), .B1(\mreg/_04751_ ), .B2(\mreg/_02817_ ), .ZN(\mreg/_03233_ ) );
NAND4_X1 \mreg/_09154_ ( .A1(\mreg/_03230_ ), .A2(\mreg/_03231_ ), .A3(\mreg/_03232_ ), .A4(\mreg/_03233_ ), .ZN(\mreg/_03234_ ) );
AND3_X1 \mreg/_09155_ ( .A1(\mreg/_02444_ ), .A2(\mreg/_04879_ ), .A3(\mreg/_02480_ ), .ZN(\mreg/_03235_ ) );
AOI21_X1 \mreg/_09156_ ( .A(\mreg/_03235_ ), .B1(\mreg/_02735_ ), .B2(\mreg/_04911_ ), .ZN(\mreg/_03236_ ) );
NAND3_X1 \mreg/_09157_ ( .A1(\mreg/_02477_ ), .A2(\mreg/_03951_ ), .A3(\mreg/_02747_ ), .ZN(\mreg/_03237_ ) );
OAI211_X2 \mreg/_09158_ ( .A(\mreg/_03236_ ), .B(\mreg/_03237_ ), .C1(\mreg/_01899_ ), .C2(\mreg/_02739_ ), .ZN(\mreg/_03238_ ) );
NAND3_X1 \mreg/_09159_ ( .A1(\mreg/_02432_ ), .A2(\mreg/_04079_ ), .A3(\mreg/_02745_ ), .ZN(\mreg/_03239_ ) );
NAND3_X1 \mreg/_09160_ ( .A1(\mreg/_02441_ ), .A2(\mreg/_04047_ ), .A3(\mreg/_02747_ ), .ZN(\mreg/_03240_ ) );
NAND3_X1 \mreg/_09161_ ( .A1(\mreg/_02426_ ), .A2(\mreg/_04111_ ), .A3(\mreg/_02747_ ), .ZN(\mreg/_03241_ ) );
NAND3_X1 \mreg/_09162_ ( .A1(\mreg/_02629_ ), .A2(\mreg/_04015_ ), .A3(\mreg/_02532_ ), .ZN(\mreg/_03242_ ) );
NAND4_X1 \mreg/_09163_ ( .A1(\mreg/_03239_ ), .A2(\mreg/_03240_ ), .A3(\mreg/_03241_ ), .A4(\mreg/_03242_ ), .ZN(\mreg/_03243_ ) );
OR4_X1 \mreg/_09164_ ( .A1(\mreg/_03228_ ), .A2(\mreg/_03234_ ), .A3(\mreg/_03238_ ), .A4(\mreg/_03243_ ), .ZN(\mreg/_03887_ ) );
NAND3_X1 \mreg/_09165_ ( .A1(\mreg/_02531_ ), .A2(\mreg/_04560_ ), .A3(\mreg/_02533_ ), .ZN(\mreg/_03244_ ) );
NAND4_X1 \mreg/_09166_ ( .A1(\mreg/_03015_ ), .A2(\mreg/_02879_ ), .A3(\mreg/_04496_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03245_ ) );
OAI21_X1 \mreg/_09167_ ( .A(\mreg/_03245_ ), .B1(\mreg/_02538_ ), .B2(\mreg/_01937_ ), .ZN(\mreg/_03246_ ) );
AOI221_X4 \mreg/_09168_ ( .A(\mreg/_03246_ ), .B1(\mreg/_04464_ ), .B2(\mreg/_02759_ ), .C1(\mreg/_04432_ ), .C2(\mreg/_02760_ ), .ZN(\mreg/_03247_ ) );
NAND3_X1 \mreg/_09169_ ( .A1(\mreg/_02546_ ), .A2(\mreg/_04592_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03248_ ) );
AND3_X1 \mreg/_09170_ ( .A1(\mreg/_02571_ ), .A2(\mreg/_04656_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03249_ ) );
AOI21_X1 \mreg/_09171_ ( .A(\mreg/_03249_ ), .B1(\mreg/_01934_ ), .B2(\mreg/_02550_ ), .ZN(\mreg/_03250_ ) );
AND4_X1 \mreg/_09172_ ( .A1(\mreg/_03244_ ), .A2(\mreg/_03247_ ), .A3(\mreg/_03248_ ), .A4(\mreg/_03250_ ), .ZN(\mreg/_03251_ ) );
NAND3_X1 \mreg/_09173_ ( .A1(\mreg/_02672_ ), .A2(\mreg/_04368_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03252_ ) );
NAND4_X1 \mreg/_09174_ ( .A1(\mreg/_02608_ ), .A2(\mreg/_04208_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02499_ ), .ZN(\mreg/_03253_ ) );
OAI21_X1 \mreg/_09175_ ( .A(\mreg/_03253_ ), .B1(\mreg/_02611_ ), .B2(\mreg/_01945_ ), .ZN(\mreg/_03254_ ) );
AOI221_X1 \mreg/_09176_ ( .A(\mreg/_03254_ ), .B1(\mreg/_04176_ ), .B2(\mreg/_02613_ ), .C1(\mreg/_04144_ ), .C2(\mreg/_02500_ ), .ZN(\mreg/_03255_ ) );
NAND3_X1 \mreg/_09177_ ( .A1(\mreg/_02674_ ), .A2(\mreg/_04400_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03256_ ) );
AND3_X1 \mreg/_09178_ ( .A1(\mreg/_02520_ ), .A2(\mreg/_04304_ ), .A3(\mreg/_02568_ ), .ZN(\mreg/_03257_ ) );
AOI21_X1 \mreg/_09179_ ( .A(\mreg/_03257_ ), .B1(\mreg/_04336_ ), .B2(\mreg/_02947_ ), .ZN(\mreg/_03258_ ) );
AND4_X1 \mreg/_09180_ ( .A1(\mreg/_03252_ ), .A2(\mreg/_03255_ ), .A3(\mreg/_03256_ ), .A4(\mreg/_03258_ ), .ZN(\mreg/_03259_ ) );
NAND3_X1 \mreg/_09181_ ( .A1(\mreg/_02583_ ), .A2(\mreg/_04272_ ), .A3(\mreg/_02820_ ), .ZN(\mreg/_03260_ ) );
AND3_X1 \mreg/_09182_ ( .A1(\mreg/_02632_ ), .A2(\mreg/_04848_ ), .A3(\mreg/_02566_ ), .ZN(\mreg/_03261_ ) );
AOI21_X1 \mreg/_09183_ ( .A(\mreg/_03261_ ), .B1(\mreg/_04816_ ), .B2(\mreg/_02636_ ), .ZN(\mreg/_03262_ ) );
AOI22_X1 \mreg/_09184_ ( .A1(\mreg/_04624_ ), .A2(\mreg/_02724_ ), .B1(\mreg/_02723_ ), .B2(\mreg/_04720_ ), .ZN(\mreg/_03263_ ) );
AOI22_X1 \mreg/_09185_ ( .A1(\mreg/_02815_ ), .A2(\mreg/_04784_ ), .B1(\mreg/_04752_ ), .B2(\mreg/_02817_ ), .ZN(\mreg/_03264_ ) );
AND4_X1 \mreg/_09186_ ( .A1(\mreg/_03260_ ), .A2(\mreg/_03262_ ), .A3(\mreg/_03263_ ), .A4(\mreg/_03264_ ), .ZN(\mreg/_03265_ ) );
NAND3_X1 \mreg/_09187_ ( .A1(\mreg/_02641_ ), .A2(\mreg/_03952_ ), .A3(\mreg/_02642_ ), .ZN(\mreg/_03266_ ) );
NAND3_X1 \mreg/_09188_ ( .A1(\mreg/_02629_ ), .A2(\mreg/_04016_ ), .A3(\mreg/_02448_ ), .ZN(\mreg/_03267_ ) );
NAND3_X1 \mreg/_09189_ ( .A1(\mreg/_02571_ ), .A2(\mreg/_04080_ ), .A3(\mreg/_02486_ ), .ZN(\mreg/_03268_ ) );
NAND3_X1 \mreg/_09190_ ( .A1(\mreg/_02696_ ), .A2(\mreg/_04048_ ), .A3(\mreg/_02572_ ), .ZN(\mreg/_03269_ ) );
NAND3_X1 \mreg/_09191_ ( .A1(\mreg/_02699_ ), .A2(\mreg/_04112_ ), .A3(\mreg/_02633_ ), .ZN(\mreg/_03270_ ) );
AND4_X1 \mreg/_09192_ ( .A1(\mreg/_03267_ ), .A2(\mreg/_03268_ ), .A3(\mreg/_03269_ ), .A4(\mreg/_03270_ ), .ZN(\mreg/_03271_ ) );
NAND3_X1 \mreg/_09193_ ( .A1(\mreg/_02647_ ), .A2(\mreg/_03984_ ), .A3(\mreg/_02654_ ), .ZN(\mreg/_03272_ ) );
AND3_X1 \mreg/_09194_ ( .A1(\mreg/_02729_ ), .A2(\mreg/_04880_ ), .A3(\mreg/_02644_ ), .ZN(\mreg/_03273_ ) );
AOI21_X1 \mreg/_09195_ ( .A(\mreg/_03273_ ), .B1(\mreg/_02735_ ), .B2(\mreg/_04912_ ), .ZN(\mreg/_03274_ ) );
AND4_X1 \mreg/_09196_ ( .A1(\mreg/_03266_ ), .A2(\mreg/_03271_ ), .A3(\mreg/_03272_ ), .A4(\mreg/_03274_ ), .ZN(\mreg/_03275_ ) );
NAND4_X1 \mreg/_09197_ ( .A1(\mreg/_03251_ ), .A2(\mreg/_03259_ ), .A3(\mreg/_03265_ ), .A4(\mreg/_03275_ ), .ZN(\mreg/_03888_ ) );
NAND3_X1 \mreg/_09198_ ( .A1(\mreg/_02597_ ), .A2(\mreg/_04594_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03276_ ) );
NAND3_X1 \mreg/_09199_ ( .A1(\mreg/_02599_ ), .A2(\mreg/_04562_ ), .A3(\mreg/_02446_ ), .ZN(\mreg/_03277_ ) );
NAND2_X1 \mreg/_09200_ ( .A1(\mreg/_03276_ ), .A2(\mreg/_03277_ ), .ZN(\mreg/_03278_ ) );
AOI221_X4 \mreg/_09201_ ( .A(\mreg/_03278_ ), .B1(\mreg/_01970_ ), .B2(\mreg/_02549_ ), .C1(\mreg/_04658_ ), .C2(\mreg/_02603_ ), .ZN(\mreg/_03279_ ) );
NAND4_X1 \mreg/_09202_ ( .A1(\mreg/_03015_ ), .A2(\mreg/_02879_ ), .A3(\mreg/_04498_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03280_ ) );
OAI21_X1 \mreg/_09203_ ( .A(\mreg/_03280_ ), .B1(\mreg/_02538_ ), .B2(\mreg/_01974_ ), .ZN(\mreg/_03281_ ) );
AOI221_X4 \mreg/_09204_ ( .A(\mreg/_03281_ ), .B1(\mreg/_04466_ ), .B2(\mreg/_02759_ ), .C1(\mreg/_04434_ ), .C2(\mreg/_02760_ ), .ZN(\mreg/_03282_ ) );
NAND4_X1 \mreg/_09205_ ( .A1(\mreg/_02585_ ), .A2(\mreg/_04210_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02609_ ), .ZN(\mreg/_03283_ ) );
NAND4_X1 \mreg/_09206_ ( .A1(\mreg/_02413_ ), .A2(\mreg/_02579_ ), .A3(\mreg/_04242_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03284_ ) );
NAND2_X1 \mreg/_09207_ ( .A1(\mreg/_03283_ ), .A2(\mreg/_03284_ ), .ZN(\mreg/_03285_ ) );
AOI221_X4 \mreg/_09208_ ( .A(\mreg/_03285_ ), .B1(\mreg/_04178_ ), .B2(\mreg/_02613_ ), .C1(\mreg/_04146_ ), .C2(\mreg/_02614_ ), .ZN(\mreg/_03286_ ) );
NAND3_X1 \mreg/_09209_ ( .A1(\mreg/_02715_ ), .A2(\mreg/_04370_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03287_ ) );
NAND3_X1 \mreg/_09210_ ( .A1(\mreg/_02565_ ), .A2(\mreg/_04402_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03288_ ) );
NAND3_X1 \mreg/_09211_ ( .A1(\mreg/_02767_ ), .A2(\mreg/_04338_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03289_ ) );
NAND3_X1 \mreg/_09212_ ( .A1(\mreg/_02520_ ), .A2(\mreg/_04306_ ), .A3(\mreg/_02467_ ), .ZN(\mreg/_03290_ ) );
AND4_X1 \mreg/_09213_ ( .A1(\mreg/_03287_ ), .A2(\mreg/_03288_ ), .A3(\mreg/_03289_ ), .A4(\mreg/_03290_ ), .ZN(\mreg/_03291_ ) );
AND4_X1 \mreg/_09214_ ( .A1(\mreg/_03279_ ), .A2(\mreg/_03282_ ), .A3(\mreg/_03286_ ), .A4(\mreg/_03291_ ), .ZN(\mreg/_03292_ ) );
NAND3_X1 \mreg/_09215_ ( .A1(\mreg/_02455_ ), .A2(\mreg/_04818_ ), .A3(\mreg/_02779_ ), .ZN(\mreg/_03293_ ) );
NAND3_X1 \mreg/_09216_ ( .A1(\mreg/_02842_ ), .A2(\mreg/_04850_ ), .A3(\mreg/_02779_ ), .ZN(\mreg/_03294_ ) );
NAND3_X1 \mreg/_09217_ ( .A1(\mreg/_02503_ ), .A2(\mreg/_04786_ ), .A3(\mreg/_02779_ ), .ZN(\mreg/_03295_ ) );
NAND3_X1 \mreg/_09218_ ( .A1(\mreg/_02730_ ), .A2(\mreg/_02512_ ), .A3(\mreg/_04754_ ), .ZN(\mreg/_03296_ ) );
NAND4_X1 \mreg/_09219_ ( .A1(\mreg/_03293_ ), .A2(\mreg/_03294_ ), .A3(\mreg/_03295_ ), .A4(\mreg/_03296_ ), .ZN(\mreg/_03297_ ) );
AND3_X1 \mreg/_09220_ ( .A1(\mreg/_02845_ ), .A2(\mreg/_04274_ ), .A3(\mreg/_02737_ ), .ZN(\mreg/_03298_ ) );
AND3_X1 \mreg/_09221_ ( .A1(\mreg/_02490_ ), .A2(\mreg/_04626_ ), .A3(\mreg/_02737_ ), .ZN(\mreg/_03299_ ) );
AND3_X1 \mreg/_09222_ ( .A1(\mreg/_02855_ ), .A2(\mreg/_04722_ ), .A3(\mreg/_02745_ ), .ZN(\mreg/_03300_ ) );
NOR4_X1 \mreg/_09223_ ( .A1(\mreg/_03297_ ), .A2(\mreg/_03298_ ), .A3(\mreg/_03299_ ), .A4(\mreg/_03300_ ), .ZN(\mreg/_03301_ ) );
NAND3_X1 \mreg/_09224_ ( .A1(\mreg/_02639_ ), .A2(\mreg/_04914_ ), .A3(\mreg/_02820_ ), .ZN(\mreg/_03302_ ) );
NAND3_X1 \mreg/_09225_ ( .A1(\mreg/_02641_ ), .A2(\mreg/_03954_ ), .A3(\mreg/_02642_ ), .ZN(\mreg/_03303_ ) );
NAND3_X1 \mreg/_09226_ ( .A1(\mreg/_02630_ ), .A2(\mreg/_02645_ ), .A3(\mreg/_04882_ ), .ZN(\mreg/_03304_ ) );
NAND3_X1 \mreg/_09227_ ( .A1(\mreg/_02647_ ), .A2(\mreg/_03986_ ), .A3(\mreg/_02648_ ), .ZN(\mreg/_03305_ ) );
AND4_X1 \mreg/_09228_ ( .A1(\mreg/_03302_ ), .A2(\mreg/_03303_ ), .A3(\mreg/_03304_ ), .A4(\mreg/_03305_ ), .ZN(\mreg/_03306_ ) );
NAND3_X1 \mreg/_09229_ ( .A1(\mreg/_02630_ ), .A2(\mreg/_04018_ ), .A3(\mreg/_02742_ ), .ZN(\mreg/_03307_ ) );
NAND3_X1 \mreg/_09230_ ( .A1(\mreg/_02785_ ), .A2(\mreg/_04082_ ), .A3(\mreg/_02652_ ), .ZN(\mreg/_03308_ ) );
NAND3_X1 \mreg/_09231_ ( .A1(\mreg/_02744_ ), .A2(\mreg/_04050_ ), .A3(\mreg/_02654_ ), .ZN(\mreg/_03309_ ) );
NAND3_X1 \mreg/_09232_ ( .A1(\mreg/_02787_ ), .A2(\mreg/_04114_ ), .A3(\mreg/_02779_ ), .ZN(\mreg/_03310_ ) );
AND4_X1 \mreg/_09233_ ( .A1(\mreg/_03307_ ), .A2(\mreg/_03308_ ), .A3(\mreg/_03309_ ), .A4(\mreg/_03310_ ), .ZN(\mreg/_03311_ ) );
NAND4_X1 \mreg/_09234_ ( .A1(\mreg/_03292_ ), .A2(\mreg/_03301_ ), .A3(\mreg/_03306_ ), .A4(\mreg/_03311_ ), .ZN(\mreg/_03890_ ) );
NAND3_X1 \mreg/_09235_ ( .A1(\mreg/_02516_ ), .A2(\mreg/_04659_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03312_ ) );
NAND4_X1 \mreg/_09236_ ( .A1(\mreg/_03015_ ), .A2(\mreg/_02879_ ), .A3(\mreg/_04499_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03313_ ) );
OAI21_X1 \mreg/_09237_ ( .A(\mreg/_03313_ ), .B1(\mreg/_02538_ ), .B2(\mreg/_02012_ ), .ZN(\mreg/_03314_ ) );
AOI221_X4 \mreg/_09238_ ( .A(\mreg/_03314_ ), .B1(\mreg/_04467_ ), .B2(\mreg/_02759_ ), .C1(\mreg/_04435_ ), .C2(\mreg/_02760_ ), .ZN(\mreg/_03315_ ) );
NAND3_X1 \mreg/_09239_ ( .A1(\mreg/_02524_ ), .A2(\mreg/_02008_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03316_ ) );
AND3_X1 \mreg/_09240_ ( .A1(\mreg/_02619_ ), .A2(\mreg/_04563_ ), .A3(\mreg/_02664_ ), .ZN(\mreg/_03317_ ) );
AOI21_X1 \mreg/_09241_ ( .A(\mreg/_03317_ ), .B1(\mreg/_02527_ ), .B2(\mreg/_04595_ ), .ZN(\mreg/_03318_ ) );
AND4_X1 \mreg/_09242_ ( .A1(\mreg/_03312_ ), .A2(\mreg/_03315_ ), .A3(\mreg/_03316_ ), .A4(\mreg/_03318_ ), .ZN(\mreg/_03319_ ) );
NAND4_X1 \mreg/_09243_ ( .A1(\mreg/_02586_ ), .A2(\mreg/_04211_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02579_ ), .ZN(\mreg/_03320_ ) );
NAND4_X1 \mreg/_09244_ ( .A1(\mreg/_02589_ ), .A2(\mreg/_02580_ ), .A3(\mreg/_04243_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03321_ ) );
NAND2_X1 \mreg/_09245_ ( .A1(\mreg/_03320_ ), .A2(\mreg/_03321_ ), .ZN(\mreg/_03322_ ) );
AOI221_X4 \mreg/_09246_ ( .A(\mreg/_03322_ ), .B1(\mreg/_04179_ ), .B2(\mreg/_02496_ ), .C1(\mreg/_04147_ ), .C2(\mreg/_02501_ ), .ZN(\mreg/_03323_ ) );
NAND3_X1 \mreg/_09247_ ( .A1(\mreg/_02506_ ), .A2(\mreg/_04371_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03324_ ) );
NAND3_X1 \mreg/_09248_ ( .A1(\mreg/_02674_ ), .A2(\mreg/_04403_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03325_ ) );
NAND3_X1 \mreg/_09249_ ( .A1(\mreg/_02504_ ), .A2(\mreg/_04339_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03326_ ) );
NAND3_X1 \mreg/_09250_ ( .A1(\mreg/_02511_ ), .A2(\mreg/_04307_ ), .A3(\mreg/_02513_ ), .ZN(\mreg/_03327_ ) );
AND4_X1 \mreg/_09251_ ( .A1(\mreg/_03324_ ), .A2(\mreg/_03325_ ), .A3(\mreg/_03326_ ), .A4(\mreg/_03327_ ), .ZN(\mreg/_03328_ ) );
AND3_X1 \mreg/_09252_ ( .A1(\mreg/_02855_ ), .A2(\mreg/_04723_ ), .A3(\mreg/_02415_ ), .ZN(\mreg/_03329_ ) );
AOI221_X4 \mreg/_09253_ ( .A(\mreg/_03329_ ), .B1(\mreg/_02627_ ), .B2(\mreg/_04627_ ), .C1(\mreg/_04275_ ), .C2(\mreg/_02420_ ), .ZN(\mreg/_03330_ ) );
NAND3_X1 \mreg/_09254_ ( .A1(\mreg/_02463_ ), .A2(\mreg/_04787_ ), .A3(\mreg/_02460_ ), .ZN(\mreg/_03331_ ) );
NAND3_X1 \mreg/_09255_ ( .A1(\mreg/_02454_ ), .A2(\mreg/_04819_ ), .A3(\mreg/_02486_ ), .ZN(\mreg/_03332_ ) );
NAND3_X1 \mreg/_09256_ ( .A1(\mreg/_02632_ ), .A2(\mreg/_04851_ ), .A3(\mreg/_02572_ ), .ZN(\mreg/_03333_ ) );
NAND3_X1 \mreg/_09257_ ( .A1(\mreg/_02684_ ), .A2(\mreg/_02568_ ), .A3(\mreg/_04755_ ), .ZN(\mreg/_03334_ ) );
AND4_X1 \mreg/_09258_ ( .A1(\mreg/_03331_ ), .A2(\mreg/_03332_ ), .A3(\mreg/_03333_ ), .A4(\mreg/_03334_ ), .ZN(\mreg/_03335_ ) );
NAND3_X1 \mreg/_09259_ ( .A1(\mreg/_02471_ ), .A2(\mreg/_04915_ ), .A3(\mreg/_02464_ ), .ZN(\mreg/_03336_ ) );
NAND3_X1 \mreg/_09260_ ( .A1(\mreg/_02476_ ), .A2(\mreg/_03955_ ), .A3(\mreg/_02688_ ), .ZN(\mreg/_03337_ ) );
NAND3_X1 \mreg/_09261_ ( .A1(\mreg/_02729_ ), .A2(\mreg/_02644_ ), .A3(\mreg/_04883_ ), .ZN(\mreg/_03338_ ) );
NAND3_X1 \mreg/_09262_ ( .A1(\mreg/_02484_ ), .A2(\mreg/_03987_ ), .A3(\mreg/_02691_ ), .ZN(\mreg/_03339_ ) );
AND4_X1 \mreg/_09263_ ( .A1(\mreg/_03336_ ), .A2(\mreg/_03337_ ), .A3(\mreg/_03338_ ), .A4(\mreg/_03339_ ), .ZN(\mreg/_03340_ ) );
NAND3_X1 \mreg/_09264_ ( .A1(\mreg/_02479_ ), .A2(\mreg/_04019_ ), .A3(\mreg/_02664_ ), .ZN(\mreg/_03341_ ) );
NAND3_X1 \mreg/_09265_ ( .A1(\mreg/_02431_ ), .A2(\mreg/_04083_ ), .A3(\mreg/_02691_ ), .ZN(\mreg/_03342_ ) );
NAND3_X1 \mreg/_09266_ ( .A1(\mreg/_02440_ ), .A2(\mreg/_04051_ ), .A3(\mreg/_02697_ ), .ZN(\mreg/_03343_ ) );
NAND3_X1 \mreg/_09267_ ( .A1(\mreg/_02425_ ), .A2(\mreg/_04115_ ), .A3(\mreg/_02700_ ), .ZN(\mreg/_03344_ ) );
AND4_X1 \mreg/_09268_ ( .A1(\mreg/_03341_ ), .A2(\mreg/_03342_ ), .A3(\mreg/_03343_ ), .A4(\mreg/_03344_ ), .ZN(\mreg/_03345_ ) );
AND4_X2 \mreg/_09269_ ( .A1(\mreg/_03330_ ), .A2(\mreg/_03335_ ), .A3(\mreg/_03340_ ), .A4(\mreg/_03345_ ), .ZN(\mreg/_03346_ ) );
NAND4_X1 \mreg/_09270_ ( .A1(\mreg/_03319_ ), .A2(\mreg/_03323_ ), .A3(\mreg/_03328_ ), .A4(\mreg/_03346_ ), .ZN(\mreg/_03891_ ) );
AND3_X1 \mreg/_09271_ ( .A1(\mreg/_02855_ ), .A2(\mreg/_04724_ ), .A3(\mreg/_02411_ ), .ZN(\mreg/_03347_ ) );
AOI221_X1 \mreg/_09272_ ( .A(\mreg/_03347_ ), .B1(\mreg/_02724_ ), .B2(\mreg/_04628_ ), .C1(\mreg/_04276_ ), .C2(\mreg/_02421_ ), .ZN(\mreg/_03348_ ) );
NAND3_X1 \mreg/_09273_ ( .A1(\mreg/_02453_ ), .A2(\mreg/_04820_ ), .A3(\mreg/_02411_ ), .ZN(\mreg/_03349_ ) );
NAND3_X1 \mreg/_09274_ ( .A1(\mreg/_02458_ ), .A2(\mreg/_04852_ ), .A3(\mreg/_02553_ ), .ZN(\mreg/_03350_ ) );
NAND2_X1 \mreg/_09275_ ( .A1(\mreg/_03349_ ), .A2(\mreg/_03350_ ), .ZN(\mreg/_03351_ ) );
AOI221_X4 \mreg/_09276_ ( .A(\mreg/_03351_ ), .B1(\mreg/_04788_ ), .B2(\mreg/_02814_ ), .C1(\mreg/_04756_ ), .C2(\mreg/_02817_ ), .ZN(\mreg/_03352_ ) );
NAND3_X1 \mreg/_09277_ ( .A1(\mreg/_02472_ ), .A2(\mreg/_04916_ ), .A3(\mreg/_02428_ ), .ZN(\mreg/_03353_ ) );
NAND3_X1 \mreg/_09278_ ( .A1(\mreg/_02477_ ), .A2(\mreg/_03956_ ), .A3(\mreg/_02460_ ), .ZN(\mreg/_03354_ ) );
NAND3_X1 \mreg/_09279_ ( .A1(\mreg/_02445_ ), .A2(\mreg/_02851_ ), .A3(\mreg/_04884_ ), .ZN(\mreg/_03355_ ) );
NAND3_X1 \mreg/_09280_ ( .A1(\mreg/_02485_ ), .A2(\mreg/_03988_ ), .A3(\mreg/_02563_ ), .ZN(\mreg/_03356_ ) );
AND4_X1 \mreg/_09281_ ( .A1(\mreg/_03353_ ), .A2(\mreg/_03354_ ), .A3(\mreg/_03355_ ), .A4(\mreg/_03356_ ), .ZN(\mreg/_03357_ ) );
NAND3_X1 \mreg/_09282_ ( .A1(\mreg/_02629_ ), .A2(\mreg/_04020_ ), .A3(\mreg/_02448_ ), .ZN(\mreg/_03358_ ) );
NAND3_X1 \mreg/_09283_ ( .A1(\mreg/_02432_ ), .A2(\mreg/_04084_ ), .A3(\mreg/_02464_ ), .ZN(\mreg/_03359_ ) );
NAND3_X1 \mreg/_09284_ ( .A1(\mreg/_02441_ ), .A2(\mreg/_04052_ ), .A3(\mreg/_02563_ ), .ZN(\mreg/_03360_ ) );
NAND3_X1 \mreg/_09285_ ( .A1(\mreg/_02699_ ), .A2(\mreg/_04116_ ), .A3(\mreg/_02486_ ), .ZN(\mreg/_03361_ ) );
AND4_X1 \mreg/_09286_ ( .A1(\mreg/_03358_ ), .A2(\mreg/_03359_ ), .A3(\mreg/_03360_ ), .A4(\mreg/_03361_ ), .ZN(\mreg/_03362_ ) );
AND4_X1 \mreg/_09287_ ( .A1(\mreg/_03348_ ), .A2(\mreg/_03352_ ), .A3(\mreg/_03357_ ), .A4(\mreg/_03362_ ), .ZN(\mreg/_03363_ ) );
NAND3_X1 \mreg/_09288_ ( .A1(\mreg/_02531_ ), .A2(\mreg/_04564_ ), .A3(\mreg/_02533_ ), .ZN(\mreg/_03364_ ) );
NAND3_X1 \mreg/_09289_ ( .A1(\mreg/_02516_ ), .A2(\mreg/_04660_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03365_ ) );
NAND3_X1 \mreg/_09290_ ( .A1(\mreg/_02546_ ), .A2(\mreg/_04596_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03366_ ) );
NAND3_X1 \mreg/_09291_ ( .A1(\mreg/_02524_ ), .A2(\mreg/_02043_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03367_ ) );
AND4_X1 \mreg/_09292_ ( .A1(\mreg/_03364_ ), .A2(\mreg/_03365_ ), .A3(\mreg/_03366_ ), .A4(\mreg/_03367_ ), .ZN(\mreg/_03368_ ) );
NAND4_X1 \mreg/_09293_ ( .A1(\mreg/_02585_ ), .A2(\mreg/_02644_ ), .A3(\mreg/_04500_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03369_ ) );
OAI21_X1 \mreg/_09294_ ( .A(\mreg/_03369_ ), .B1(\mreg/_02539_ ), .B2(\mreg/_02047_ ), .ZN(\mreg/_03370_ ) );
AOI221_X4 \mreg/_09295_ ( .A(\mreg/_03370_ ), .B1(\mreg/_04468_ ), .B2(\mreg/_02542_ ), .C1(\mreg/_04436_ ), .C2(\mreg/_02544_ ), .ZN(\mreg/_03371_ ) );
NAND3_X1 \mreg/_09296_ ( .A1(\mreg/_02506_ ), .A2(\mreg/_04372_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03372_ ) );
NAND4_X1 \mreg/_09297_ ( .A1(\mreg/_02585_ ), .A2(\mreg/_04212_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02609_ ), .ZN(\mreg/_03373_ ) );
NAND4_X1 \mreg/_09298_ ( .A1(\mreg/_02413_ ), .A2(\mreg/_02609_ ), .A3(\mreg/_04244_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03374_ ) );
NAND2_X1 \mreg/_09299_ ( .A1(\mreg/_03373_ ), .A2(\mreg/_03374_ ), .ZN(\mreg/_03375_ ) );
AOI221_X4 \mreg/_09300_ ( .A(\mreg/_03375_ ), .B1(\mreg/_04180_ ), .B2(\mreg/_02495_ ), .C1(\mreg/_04148_ ), .C2(\mreg/_02500_ ), .ZN(\mreg/_03376_ ) );
NAND3_X1 \mreg/_09301_ ( .A1(\mreg/_02508_ ), .A2(\mreg/_04404_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03377_ ) );
AND3_X1 \mreg/_09302_ ( .A1(\mreg/_02510_ ), .A2(\mreg/_04308_ ), .A3(\mreg/_02466_ ), .ZN(\mreg/_03378_ ) );
AOI21_X1 \mreg/_09303_ ( .A(\mreg/_03378_ ), .B1(\mreg/_04340_ ), .B2(\mreg/_02947_ ), .ZN(\mreg/_03379_ ) );
AND4_X1 \mreg/_09304_ ( .A1(\mreg/_03372_ ), .A2(\mreg/_03376_ ), .A3(\mreg/_03377_ ), .A4(\mreg/_03379_ ), .ZN(\mreg/_03380_ ) );
NAND4_X1 \mreg/_09305_ ( .A1(\mreg/_03363_ ), .A2(\mreg/_03368_ ), .A3(\mreg/_03371_ ), .A4(\mreg/_03380_ ), .ZN(\mreg/_03892_ ) );
NAND3_X1 \mreg/_09306_ ( .A1(\mreg/_02639_ ), .A2(\mreg/_04469_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03381_ ) );
NAND3_X1 \mreg/_09307_ ( .A1(\mreg/_02530_ ), .A2(\mreg/_04565_ ), .A3(\mreg/_02532_ ), .ZN(\mreg/_03382_ ) );
NAND3_X1 \mreg/_09308_ ( .A1(\mreg/_02715_ ), .A2(\mreg/_04373_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03383_ ) );
NAND3_X1 \mreg/_09309_ ( .A1(\mreg/_02490_ ), .A2(\mreg/_04629_ ), .A3(\mreg/_02434_ ), .ZN(\mreg/_03384_ ) );
NAND3_X1 \mreg/_09310_ ( .A1(\mreg/_02445_ ), .A2(\mreg/_04021_ ), .A3(\mreg/_02448_ ), .ZN(\mreg/_03385_ ) );
AND4_X1 \mreg/_09311_ ( .A1(\mreg/_03382_ ), .A2(\mreg/_03383_ ), .A3(\mreg/_03384_ ), .A4(\mreg/_03385_ ), .ZN(\mreg/_03386_ ) );
NAND3_X1 \mreg/_09312_ ( .A1(\mreg/_02583_ ), .A2(\mreg/_04277_ ), .A3(\mreg/_02820_ ), .ZN(\mreg/_03387_ ) );
AOI22_X1 \mreg/_09313_ ( .A1(\mreg/_02815_ ), .A2(\mreg/_04789_ ), .B1(\mreg/_02501_ ), .B2(\mreg/_04149_ ), .ZN(\mreg/_03388_ ) );
AND4_X1 \mreg/_09314_ ( .A1(\mreg/_03381_ ), .A2(\mreg/_03386_ ), .A3(\mreg/_03387_ ), .A4(\mreg/_03388_ ), .ZN(\mreg/_03389_ ) );
NAND3_X1 \mreg/_09315_ ( .A1(\mreg/_02504_ ), .A2(\mreg/_04341_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03390_ ) );
AOI22_X1 \mreg/_09316_ ( .A1(\mreg/_04821_ ), .A2(\mreg/_02636_ ), .B1(\mreg/_02735_ ), .B2(\mreg/_04917_ ), .ZN(\mreg/_03391_ ) );
AOI22_X1 \mreg/_09317_ ( .A1(\mreg/_02603_ ), .A2(\mreg/_04661_ ), .B1(\mreg/_02807_ ), .B2(\mreg/_04309_ ), .ZN(\mreg/_03392_ ) );
AOI22_X1 \mreg/_09318_ ( .A1(\mreg/_02560_ ), .A2(\mreg/_03957_ ), .B1(\mreg/_02550_ ), .B2(\mreg/_02089_ ), .ZN(\mreg/_03393_ ) );
AND4_X1 \mreg/_09319_ ( .A1(\mreg/_03390_ ), .A2(\mreg/_03391_ ), .A3(\mreg/_03392_ ), .A4(\mreg/_03393_ ), .ZN(\mreg/_03394_ ) );
NAND3_X1 \mreg/_09320_ ( .A1(\mreg/_02730_ ), .A2(\mreg/_02512_ ), .A3(\mreg/_04757_ ), .ZN(\mreg/_03395_ ) );
OAI21_X1 \mreg/_09321_ ( .A(\mreg/_03395_ ), .B1(\mreg/_03112_ ), .B2(\mreg/_02079_ ), .ZN(\mreg/_03396_ ) );
NAND4_X1 \mreg/_09322_ ( .A1(\mreg/_02587_ ), .A2(\mreg/_02838_ ), .A3(\mreg/_04501_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03397_ ) );
OAI21_X1 \mreg/_09323_ ( .A(\mreg/_03397_ ), .B1(\mreg/_02539_ ), .B2(\mreg/_02087_ ), .ZN(\mreg/_03398_ ) );
NAND4_X1 \mreg/_09324_ ( .A1(\mreg/_02587_ ), .A2(\mreg/_04213_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02580_ ), .ZN(\mreg/_03399_ ) );
OAI21_X1 \mreg/_09325_ ( .A(\mreg/_03399_ ), .B1(\mreg/_02493_ ), .B2(\mreg/_02092_ ), .ZN(\mreg/_03400_ ) );
NAND3_X1 \mreg/_09326_ ( .A1(\mreg/_02787_ ), .A2(\mreg/_04117_ ), .A3(\mreg/_02747_ ), .ZN(\mreg/_03401_ ) );
OAI21_X1 \mreg/_09327_ ( .A(\mreg/_03401_ ), .B1(\mreg/_03116_ ), .B2(\mreg/_02083_ ), .ZN(\mreg/_03402_ ) );
NOR4_X1 \mreg/_09328_ ( .A1(\mreg/_03396_ ), .A2(\mreg/_03398_ ), .A3(\mreg/_03400_ ), .A4(\mreg/_03402_ ), .ZN(\mreg/_03403_ ) );
OAI22_X1 \mreg/_09329_ ( .A1(\mreg/_02102_ ), .A2(\mreg/_02749_ ), .B1(\mreg/_02739_ ), .B2(\mreg/_02103_ ), .ZN(\mreg/_03404_ ) );
NAND3_X1 \mreg/_09330_ ( .A1(\mreg/_02842_ ), .A2(\mreg/_04405_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03405_ ) );
NAND3_X1 \mreg/_09331_ ( .A1(\mreg/_02441_ ), .A2(\mreg/_04597_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03406_ ) );
NAND3_X1 \mreg/_09332_ ( .A1(\mreg/_02837_ ), .A2(\mreg/_04437_ ), .A3(\mreg/_02838_ ), .ZN(\mreg/_03407_ ) );
NAND3_X1 \mreg/_09333_ ( .A1(\mreg/_02845_ ), .A2(\mreg/_04181_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03408_ ) );
NAND4_X1 \mreg/_09334_ ( .A1(\mreg/_03405_ ), .A2(\mreg/_03406_ ), .A3(\mreg/_03407_ ), .A4(\mreg/_03408_ ), .ZN(\mreg/_03409_ ) );
AND3_X1 \mreg/_09335_ ( .A1(\mreg/_02842_ ), .A2(\mreg/_04853_ ), .A3(\mreg/_02745_ ), .ZN(\mreg/_03410_ ) );
AND3_X1 \mreg/_09336_ ( .A1(\mreg/_02741_ ), .A2(\mreg/_04885_ ), .A3(\mreg/_02838_ ), .ZN(\mreg/_03411_ ) );
NOR4_X1 \mreg/_09337_ ( .A1(\mreg/_03404_ ), .A2(\mreg/_03409_ ), .A3(\mreg/_03410_ ), .A4(\mreg/_03411_ ), .ZN(\mreg/_03412_ ) );
NAND4_X1 \mreg/_09338_ ( .A1(\mreg/_03389_ ), .A2(\mreg/_03394_ ), .A3(\mreg/_03403_ ), .A4(\mreg/_03412_ ), .ZN(\mreg/_03893_ ) );
NAND3_X1 \mreg/_09339_ ( .A1(\mreg/_02672_ ), .A2(\mreg/_04374_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03413_ ) );
NAND4_X1 \mreg/_09340_ ( .A1(\mreg/_02585_ ), .A2(\mreg/_04214_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02579_ ), .ZN(\mreg/_03414_ ) );
NAND4_X1 \mreg/_09341_ ( .A1(\mreg/_02413_ ), .A2(\mreg/_02579_ ), .A3(\mreg/_04246_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03415_ ) );
NAND2_X1 \mreg/_09342_ ( .A1(\mreg/_03414_ ), .A2(\mreg/_03415_ ), .ZN(\mreg/_03416_ ) );
AOI221_X4 \mreg/_09343_ ( .A(\mreg/_03416_ ), .B1(\mreg/_04182_ ), .B2(\mreg/_02496_ ), .C1(\mreg/_04150_ ), .C2(\mreg/_02501_ ), .ZN(\mreg/_03417_ ) );
NAND3_X1 \mreg/_09344_ ( .A1(\mreg/_02674_ ), .A2(\mreg/_04406_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03418_ ) );
AND3_X1 \mreg/_09345_ ( .A1(\mreg/_02767_ ), .A2(\mreg/_04342_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03419_ ) );
AOI21_X1 \mreg/_09346_ ( .A(\mreg/_03419_ ), .B1(\mreg/_04310_ ), .B2(\mreg/_02807_ ), .ZN(\mreg/_03420_ ) );
AND4_X1 \mreg/_09347_ ( .A1(\mreg/_03413_ ), .A2(\mreg/_03417_ ), .A3(\mreg/_03418_ ), .A4(\mreg/_03420_ ), .ZN(\mreg/_03421_ ) );
NAND3_X1 \mreg/_09348_ ( .A1(\mreg/_02531_ ), .A2(\mreg/_04566_ ), .A3(\mreg/_02533_ ), .ZN(\mreg/_03422_ ) );
NAND3_X1 \mreg/_09349_ ( .A1(\mreg/_02516_ ), .A2(\mreg/_04662_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03423_ ) );
NAND3_X1 \mreg/_09350_ ( .A1(\mreg/_02546_ ), .A2(\mreg/_04598_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03424_ ) );
NAND3_X1 \mreg/_09351_ ( .A1(\mreg/_02524_ ), .A2(\mreg/_02118_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03425_ ) );
AND4_X1 \mreg/_09352_ ( .A1(\mreg/_03422_ ), .A2(\mreg/_03423_ ), .A3(\mreg/_03424_ ), .A4(\mreg/_03425_ ), .ZN(\mreg/_03426_ ) );
AND3_X1 \mreg/_09353_ ( .A1(\mreg/_02855_ ), .A2(\mreg/_04726_ ), .A3(\mreg/_02553_ ), .ZN(\mreg/_03427_ ) );
AOI221_X2 \mreg/_09354_ ( .A(\mreg/_03427_ ), .B1(\mreg/_02627_ ), .B2(\mreg/_04630_ ), .C1(\mreg/_04278_ ), .C2(\mreg/_02421_ ), .ZN(\mreg/_03428_ ) );
NAND3_X1 \mreg/_09355_ ( .A1(\mreg/_02503_ ), .A2(\mreg/_04790_ ), .A3(\mreg/_02434_ ), .ZN(\mreg/_03429_ ) );
NAND3_X1 \mreg/_09356_ ( .A1(\mreg/_02715_ ), .A2(\mreg/_04822_ ), .A3(\mreg/_02563_ ), .ZN(\mreg/_03430_ ) );
NAND3_X1 \mreg/_09357_ ( .A1(\mreg/_02565_ ), .A2(\mreg/_04854_ ), .A3(\mreg/_02566_ ), .ZN(\mreg/_03431_ ) );
NAND3_X1 \mreg/_09358_ ( .A1(\mreg/_02479_ ), .A2(\mreg/_02568_ ), .A3(\mreg/_04758_ ), .ZN(\mreg/_03432_ ) );
AND4_X1 \mreg/_09359_ ( .A1(\mreg/_03429_ ), .A2(\mreg/_03430_ ), .A3(\mreg/_03431_ ), .A4(\mreg/_03432_ ), .ZN(\mreg/_03433_ ) );
NAND3_X1 \mreg/_09360_ ( .A1(\mreg/_02471_ ), .A2(\mreg/_04918_ ), .A3(\mreg/_02464_ ), .ZN(\mreg/_03434_ ) );
NAND3_X1 \mreg/_09361_ ( .A1(\mreg/_02476_ ), .A2(\mreg/_03958_ ), .A3(\mreg/_02566_ ), .ZN(\mreg/_03435_ ) );
NAND3_X1 \mreg/_09362_ ( .A1(\mreg/_02684_ ), .A2(\mreg/_02481_ ), .A3(\mreg/_04886_ ), .ZN(\mreg/_03436_ ) );
NAND3_X1 \mreg/_09363_ ( .A1(\mreg/_02485_ ), .A2(\mreg/_03990_ ), .A3(\mreg/_02691_ ), .ZN(\mreg/_03437_ ) );
AND4_X1 \mreg/_09364_ ( .A1(\mreg/_03434_ ), .A2(\mreg/_03435_ ), .A3(\mreg/_03436_ ), .A4(\mreg/_03437_ ), .ZN(\mreg/_03438_ ) );
NAND3_X1 \mreg/_09365_ ( .A1(\mreg/_02445_ ), .A2(\mreg/_04022_ ), .A3(\mreg/_02664_ ), .ZN(\mreg/_03439_ ) );
NAND3_X1 \mreg/_09366_ ( .A1(\mreg/_02571_ ), .A2(\mreg/_04086_ ), .A3(\mreg/_02688_ ), .ZN(\mreg/_03440_ ) );
NAND3_X1 \mreg/_09367_ ( .A1(\mreg/_02696_ ), .A2(\mreg/_04054_ ), .A3(\mreg/_02691_ ), .ZN(\mreg/_03441_ ) );
NAND3_X1 \mreg/_09368_ ( .A1(\mreg/_02699_ ), .A2(\mreg/_04118_ ), .A3(\mreg/_02700_ ), .ZN(\mreg/_03442_ ) );
AND4_X1 \mreg/_09369_ ( .A1(\mreg/_03439_ ), .A2(\mreg/_03440_ ), .A3(\mreg/_03441_ ), .A4(\mreg/_03442_ ), .ZN(\mreg/_03443_ ) );
AND4_X4 \mreg/_09370_ ( .A1(\mreg/_03428_ ), .A2(\mreg/_03433_ ), .A3(\mreg/_03438_ ), .A4(\mreg/_03443_ ), .ZN(\mreg/_03444_ ) );
NAND4_X1 \mreg/_09371_ ( .A1(\mreg/_02585_ ), .A2(\mreg/_02480_ ), .A3(\mreg/_04502_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03445_ ) );
OAI21_X1 \mreg/_09372_ ( .A(\mreg/_03445_ ), .B1(\mreg/_02539_ ), .B2(\mreg/_02121_ ), .ZN(\mreg/_03446_ ) );
AOI221_X4 \mreg/_09373_ ( .A(\mreg/_03446_ ), .B1(\mreg/_04470_ ), .B2(\mreg/_02542_ ), .C1(\mreg/_04438_ ), .C2(\mreg/_02544_ ), .ZN(\mreg/_03447_ ) );
NAND4_X1 \mreg/_09374_ ( .A1(\mreg/_03421_ ), .A2(\mreg/_03426_ ), .A3(\mreg/_03444_ ), .A4(\mreg/_03447_ ), .ZN(\mreg/_03894_ ) );
NAND3_X1 \mreg/_09375_ ( .A1(\mreg/_02530_ ), .A2(\mreg/_04567_ ), .A3(\mreg/_02532_ ), .ZN(\mreg/_03448_ ) );
NAND3_X1 \mreg/_09376_ ( .A1(\mreg/_02432_ ), .A2(\mreg/_04663_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03449_ ) );
NAND3_X1 \mreg/_09377_ ( .A1(\mreg/_02441_ ), .A2(\mreg/_04599_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03450_ ) );
NAND3_X1 \mreg/_09378_ ( .A1(\mreg/_02426_ ), .A2(\mreg/_02154_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03451_ ) );
AND4_X1 \mreg/_09379_ ( .A1(\mreg/_03448_ ), .A2(\mreg/_03449_ ), .A3(\mreg/_03450_ ), .A4(\mreg/_03451_ ), .ZN(\mreg/_03452_ ) );
NAND4_X1 \mreg/_09380_ ( .A1(\mreg/_03015_ ), .A2(\mreg/_04215_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02609_ ), .ZN(\mreg/_03453_ ) );
OAI21_X1 \mreg/_09381_ ( .A(\mreg/_03453_ ), .B1(\mreg/_02493_ ), .B2(\mreg/_02167_ ), .ZN(\mreg/_03454_ ) );
AOI221_X4 \mreg/_09382_ ( .A(\mreg/_03454_ ), .B1(\mreg/_04183_ ), .B2(\mreg/_02496_ ), .C1(\mreg/_04151_ ), .C2(\mreg/_02614_ ), .ZN(\mreg/_03455_ ) );
NAND3_X1 \mreg/_09383_ ( .A1(\mreg/_02472_ ), .A2(\mreg/_04471_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03456_ ) );
NAND3_X1 \mreg/_09384_ ( .A1(\mreg/_02530_ ), .A2(\mreg/_04439_ ), .A3(\mreg/_02851_ ), .ZN(\mreg/_03457_ ) );
NAND4_X1 \mreg/_09385_ ( .A1(\mreg/_02586_ ), .A2(\mreg/_02481_ ), .A3(\mreg/_04503_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03458_ ) );
NAND4_X1 \mreg/_09386_ ( .A1(\mreg/_02481_ ), .A2(\mreg/_04535_ ), .A3(\mreg/_02589_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03459_ ) );
AND4_X1 \mreg/_09387_ ( .A1(\mreg/_03456_ ), .A2(\mreg/_03457_ ), .A3(\mreg/_03458_ ), .A4(\mreg/_03459_ ), .ZN(\mreg/_03460_ ) );
NAND3_X1 \mreg/_09388_ ( .A1(\mreg/_02455_ ), .A2(\mreg/_04375_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03461_ ) );
NAND3_X1 \mreg/_09389_ ( .A1(\mreg/_02459_ ), .A2(\mreg/_04407_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03462_ ) );
NAND2_X1 \mreg/_09390_ ( .A1(\mreg/_03461_ ), .A2(\mreg/_03462_ ), .ZN(\mreg/_03463_ ) );
AND3_X1 \mreg/_09391_ ( .A1(\mreg/_02767_ ), .A2(\mreg/_04343_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03464_ ) );
AND3_X1 \mreg/_09392_ ( .A1(\mreg/_02520_ ), .A2(\mreg/_04311_ ), .A3(\mreg/_02568_ ), .ZN(\mreg/_03465_ ) );
NOR3_X1 \mreg/_09393_ ( .A1(\mreg/_03463_ ), .A2(\mreg/_03464_ ), .A3(\mreg/_03465_ ), .ZN(\mreg/_03466_ ) );
AND4_X1 \mreg/_09394_ ( .A1(\mreg/_03452_ ), .A2(\mreg/_03455_ ), .A3(\mreg/_03460_ ), .A4(\mreg/_03466_ ), .ZN(\mreg/_03467_ ) );
NAND3_X1 \mreg/_09395_ ( .A1(\mreg/_02672_ ), .A2(\mreg/_04823_ ), .A3(\mreg/_02624_ ), .ZN(\mreg/_03468_ ) );
AOI22_X1 \mreg/_09396_ ( .A1(\mreg/_02815_ ), .A2(\mreg/_04791_ ), .B1(\mreg/_04759_ ), .B2(\mreg/_02817_ ), .ZN(\mreg/_03469_ ) );
NAND3_X1 \mreg/_09397_ ( .A1(\mreg/_02508_ ), .A2(\mreg/_04855_ ), .A3(\mreg/_02652_ ), .ZN(\mreg/_03470_ ) );
NAND3_X1 \mreg/_09398_ ( .A1(\mreg/_02419_ ), .A2(\mreg/_04279_ ), .A3(\mreg/_02428_ ), .ZN(\mreg/_03471_ ) );
NAND3_X1 \mreg/_09399_ ( .A1(\mreg/_02490_ ), .A2(\mreg/_04631_ ), .A3(\mreg/_02428_ ), .ZN(\mreg/_03472_ ) );
NAND3_X1 \mreg/_09400_ ( .A1(\mreg/_02855_ ), .A2(\mreg/_04727_ ), .A3(\mreg/_02434_ ), .ZN(\mreg/_03473_ ) );
AND3_X1 \mreg/_09401_ ( .A1(\mreg/_03471_ ), .A2(\mreg/_03472_ ), .A3(\mreg/_03473_ ), .ZN(\mreg/_03474_ ) );
AND4_X1 \mreg/_09402_ ( .A1(\mreg/_03468_ ), .A2(\mreg/_03469_ ), .A3(\mreg/_03470_ ), .A4(\mreg/_03474_ ), .ZN(\mreg/_03475_ ) );
NAND3_X1 \mreg/_09403_ ( .A1(\mreg/_02639_ ), .A2(\mreg/_04919_ ), .A3(\mreg/_02820_ ), .ZN(\mreg/_03476_ ) );
NAND3_X1 \mreg/_09404_ ( .A1(\mreg/_02641_ ), .A2(\mreg/_03959_ ), .A3(\mreg/_02652_ ), .ZN(\mreg/_03477_ ) );
NAND3_X1 \mreg/_09405_ ( .A1(\mreg/_02730_ ), .A2(\mreg/_02645_ ), .A3(\mreg/_04887_ ), .ZN(\mreg/_03478_ ) );
NAND3_X1 \mreg/_09406_ ( .A1(\mreg/_02647_ ), .A2(\mreg/_03991_ ), .A3(\mreg/_02648_ ), .ZN(\mreg/_03479_ ) );
AND4_X1 \mreg/_09407_ ( .A1(\mreg/_03476_ ), .A2(\mreg/_03477_ ), .A3(\mreg/_03478_ ), .A4(\mreg/_03479_ ), .ZN(\mreg/_03480_ ) );
NAND3_X1 \mreg/_09408_ ( .A1(\mreg/_02630_ ), .A2(\mreg/_04023_ ), .A3(\mreg/_02742_ ), .ZN(\mreg/_03481_ ) );
NAND3_X1 \mreg/_09409_ ( .A1(\mreg/_02785_ ), .A2(\mreg/_04087_ ), .A3(\mreg/_02652_ ), .ZN(\mreg/_03482_ ) );
NAND3_X1 \mreg/_09410_ ( .A1(\mreg/_02744_ ), .A2(\mreg/_04055_ ), .A3(\mreg/_02654_ ), .ZN(\mreg/_03483_ ) );
NAND3_X1 \mreg/_09411_ ( .A1(\mreg/_02787_ ), .A2(\mreg/_04119_ ), .A3(\mreg/_02779_ ), .ZN(\mreg/_03484_ ) );
AND4_X1 \mreg/_09412_ ( .A1(\mreg/_03481_ ), .A2(\mreg/_03482_ ), .A3(\mreg/_03483_ ), .A4(\mreg/_03484_ ), .ZN(\mreg/_03485_ ) );
NAND4_X1 \mreg/_09413_ ( .A1(\mreg/_03467_ ), .A2(\mreg/_03475_ ), .A3(\mreg/_03480_ ), .A4(\mreg/_03485_ ), .ZN(\mreg/_03895_ ) );
NAND3_X1 \mreg/_09414_ ( .A1(\mreg/_02639_ ), .A2(\mreg/_04472_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03486_ ) );
NAND3_X1 \mreg/_09415_ ( .A1(\mreg/_02530_ ), .A2(\mreg/_04568_ ), .A3(\mreg/_02448_ ), .ZN(\mreg/_03487_ ) );
NAND3_X1 \mreg/_09416_ ( .A1(\mreg/_02715_ ), .A2(\mreg/_04376_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03488_ ) );
NAND3_X1 \mreg/_09417_ ( .A1(\mreg/_02490_ ), .A2(\mreg/_04632_ ), .A3(\mreg/_02434_ ), .ZN(\mreg/_03489_ ) );
NAND3_X1 \mreg/_09418_ ( .A1(\mreg/_02445_ ), .A2(\mreg/_04024_ ), .A3(\mreg/_02664_ ), .ZN(\mreg/_03490_ ) );
AND4_X1 \mreg/_09419_ ( .A1(\mreg/_03487_ ), .A2(\mreg/_03488_ ), .A3(\mreg/_03489_ ), .A4(\mreg/_03490_ ), .ZN(\mreg/_03491_ ) );
NAND3_X1 \mreg/_09420_ ( .A1(\mreg/_02583_ ), .A2(\mreg/_04280_ ), .A3(\mreg/_02820_ ), .ZN(\mreg/_03492_ ) );
AOI22_X1 \mreg/_09421_ ( .A1(\mreg/_02815_ ), .A2(\mreg/_04792_ ), .B1(\mreg/_02501_ ), .B2(\mreg/_04152_ ), .ZN(\mreg/_03493_ ) );
AND4_X1 \mreg/_09422_ ( .A1(\mreg/_03486_ ), .A2(\mreg/_03491_ ), .A3(\mreg/_03492_ ), .A4(\mreg/_03493_ ), .ZN(\mreg/_03494_ ) );
NAND3_X1 \mreg/_09423_ ( .A1(\mreg/_02504_ ), .A2(\mreg/_04344_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03495_ ) );
AOI22_X1 \mreg/_09424_ ( .A1(\mreg/_04824_ ), .A2(\mreg/_02636_ ), .B1(\mreg/_02735_ ), .B2(\mreg/_04920_ ), .ZN(\mreg/_03496_ ) );
AOI22_X1 \mreg/_09425_ ( .A1(\mreg/_02603_ ), .A2(\mreg/_04664_ ), .B1(\mreg/_02807_ ), .B2(\mreg/_04312_ ), .ZN(\mreg/_03497_ ) );
AOI22_X1 \mreg/_09426_ ( .A1(\mreg/_02560_ ), .A2(\mreg/_03960_ ), .B1(\mreg/_02550_ ), .B2(\mreg/_02199_ ), .ZN(\mreg/_03498_ ) );
AND4_X1 \mreg/_09427_ ( .A1(\mreg/_03495_ ), .A2(\mreg/_03496_ ), .A3(\mreg/_03497_ ), .A4(\mreg/_03498_ ), .ZN(\mreg/_03499_ ) );
NAND3_X1 \mreg/_09428_ ( .A1(\mreg/_02730_ ), .A2(\mreg/_02512_ ), .A3(\mreg/_04760_ ), .ZN(\mreg/_03500_ ) );
OAI21_X1 \mreg/_09429_ ( .A(\mreg/_03500_ ), .B1(\mreg/_03112_ ), .B2(\mreg/_02189_ ), .ZN(\mreg/_03501_ ) );
NAND4_X1 \mreg/_09430_ ( .A1(\mreg/_02587_ ), .A2(\mreg/_02838_ ), .A3(\mreg/_04504_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03502_ ) );
OAI21_X1 \mreg/_09431_ ( .A(\mreg/_03502_ ), .B1(\mreg/_02539_ ), .B2(\mreg/_02197_ ), .ZN(\mreg/_03503_ ) );
NAND4_X1 \mreg/_09432_ ( .A1(\mreg/_02587_ ), .A2(\mreg/_04216_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02580_ ), .ZN(\mreg/_03504_ ) );
OAI21_X1 \mreg/_09433_ ( .A(\mreg/_03504_ ), .B1(\mreg/_02493_ ), .B2(\mreg/_02202_ ), .ZN(\mreg/_03505_ ) );
NAND3_X1 \mreg/_09434_ ( .A1(\mreg/_02426_ ), .A2(\mreg/_04120_ ), .A3(\mreg/_02747_ ), .ZN(\mreg/_03506_ ) );
OAI21_X1 \mreg/_09435_ ( .A(\mreg/_03506_ ), .B1(\mreg/_03116_ ), .B2(\mreg/_02193_ ), .ZN(\mreg/_03507_ ) );
NOR4_X1 \mreg/_09436_ ( .A1(\mreg/_03501_ ), .A2(\mreg/_03503_ ), .A3(\mreg/_03505_ ), .A4(\mreg/_03507_ ), .ZN(\mreg/_03508_ ) );
OAI22_X1 \mreg/_09437_ ( .A1(\mreg/_02212_ ), .A2(\mreg/_02749_ ), .B1(\mreg/_02739_ ), .B2(\mreg/_02213_ ), .ZN(\mreg/_03509_ ) );
NAND3_X1 \mreg/_09438_ ( .A1(\mreg/_02842_ ), .A2(\mreg/_04408_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03510_ ) );
NAND3_X1 \mreg/_09439_ ( .A1(\mreg/_02441_ ), .A2(\mreg/_04600_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03511_ ) );
NAND3_X1 \mreg/_09440_ ( .A1(\mreg/_02837_ ), .A2(\mreg/_04440_ ), .A3(\mreg/_02838_ ), .ZN(\mreg/_03512_ ) );
NAND3_X1 \mreg/_09441_ ( .A1(\mreg/_02845_ ), .A2(\mreg/_04184_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03513_ ) );
NAND4_X1 \mreg/_09442_ ( .A1(\mreg/_03510_ ), .A2(\mreg/_03511_ ), .A3(\mreg/_03512_ ), .A4(\mreg/_03513_ ), .ZN(\mreg/_03514_ ) );
AND3_X1 \mreg/_09443_ ( .A1(\mreg/_02842_ ), .A2(\mreg/_04856_ ), .A3(\mreg/_02745_ ), .ZN(\mreg/_03515_ ) );
AND3_X1 \mreg/_09444_ ( .A1(\mreg/_02741_ ), .A2(\mreg/_04888_ ), .A3(\mreg/_02838_ ), .ZN(\mreg/_03516_ ) );
NOR4_X1 \mreg/_09445_ ( .A1(\mreg/_03509_ ), .A2(\mreg/_03514_ ), .A3(\mreg/_03515_ ), .A4(\mreg/_03516_ ), .ZN(\mreg/_03517_ ) );
NAND4_X1 \mreg/_09446_ ( .A1(\mreg/_03494_ ), .A2(\mreg/_03499_ ), .A3(\mreg/_03508_ ), .A4(\mreg/_03517_ ), .ZN(\mreg/_03896_ ) );
AND3_X1 \mreg/_09447_ ( .A1(\mreg/_02855_ ), .A2(\mreg/_04729_ ), .A3(\mreg/_02411_ ), .ZN(\mreg/_03518_ ) );
AOI221_X1 \mreg/_09448_ ( .A(\mreg/_03518_ ), .B1(\mreg/_02627_ ), .B2(\mreg/_04633_ ), .C1(\mreg/_04281_ ), .C2(\mreg/_02421_ ), .ZN(\mreg/_03519_ ) );
NAND3_X1 \mreg/_09449_ ( .A1(\mreg/_02503_ ), .A2(\mreg/_04793_ ), .A3(\mreg/_02428_ ), .ZN(\mreg/_03520_ ) );
NAND3_X1 \mreg/_09450_ ( .A1(\mreg/_02715_ ), .A2(\mreg/_04825_ ), .A3(\mreg/_02434_ ), .ZN(\mreg/_03521_ ) );
NAND3_X1 \mreg/_09451_ ( .A1(\mreg/_02459_ ), .A2(\mreg/_04857_ ), .A3(\mreg/_02460_ ), .ZN(\mreg/_03522_ ) );
NAND3_X1 \mreg/_09452_ ( .A1(\mreg/_02445_ ), .A2(\mreg/_02512_ ), .A3(\mreg/_04761_ ), .ZN(\mreg/_03523_ ) );
AND4_X1 \mreg/_09453_ ( .A1(\mreg/_03520_ ), .A2(\mreg/_03521_ ), .A3(\mreg/_03522_ ), .A4(\mreg/_03523_ ), .ZN(\mreg/_03524_ ) );
NAND3_X1 \mreg/_09454_ ( .A1(\mreg/_02472_ ), .A2(\mreg/_04921_ ), .A3(\mreg/_02428_ ), .ZN(\mreg/_03525_ ) );
NAND3_X1 \mreg/_09455_ ( .A1(\mreg/_02477_ ), .A2(\mreg/_03961_ ), .A3(\mreg/_02460_ ), .ZN(\mreg/_03526_ ) );
NAND3_X1 \mreg/_09456_ ( .A1(\mreg/_02445_ ), .A2(\mreg/_02481_ ), .A3(\mreg/_04889_ ), .ZN(\mreg/_03527_ ) );
NAND3_X1 \mreg/_09457_ ( .A1(\mreg/_02485_ ), .A2(\mreg/_03993_ ), .A3(\mreg/_02563_ ), .ZN(\mreg/_03528_ ) );
AND4_X1 \mreg/_09458_ ( .A1(\mreg/_03525_ ), .A2(\mreg/_03526_ ), .A3(\mreg/_03527_ ), .A4(\mreg/_03528_ ), .ZN(\mreg/_03529_ ) );
NAND3_X1 \mreg/_09459_ ( .A1(\mreg/_02629_ ), .A2(\mreg/_04025_ ), .A3(\mreg/_02448_ ), .ZN(\mreg/_03530_ ) );
NAND3_X1 \mreg/_09460_ ( .A1(\mreg/_02432_ ), .A2(\mreg/_04089_ ), .A3(\mreg/_02464_ ), .ZN(\mreg/_03531_ ) );
NAND3_X1 \mreg/_09461_ ( .A1(\mreg/_02696_ ), .A2(\mreg/_04057_ ), .A3(\mreg/_02563_ ), .ZN(\mreg/_03532_ ) );
NAND3_X1 \mreg/_09462_ ( .A1(\mreg/_02699_ ), .A2(\mreg/_04121_ ), .A3(\mreg/_02486_ ), .ZN(\mreg/_03533_ ) );
AND4_X1 \mreg/_09463_ ( .A1(\mreg/_03530_ ), .A2(\mreg/_03531_ ), .A3(\mreg/_03532_ ), .A4(\mreg/_03533_ ), .ZN(\mreg/_03534_ ) );
AND4_X1 \mreg/_09464_ ( .A1(\mreg/_03519_ ), .A2(\mreg/_03524_ ), .A3(\mreg/_03529_ ), .A4(\mreg/_03534_ ), .ZN(\mreg/_03535_ ) );
NAND3_X1 \mreg/_09465_ ( .A1(\mreg/_02696_ ), .A2(\mreg/_04601_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03536_ ) );
NAND3_X1 \mreg/_09466_ ( .A1(\mreg/_02520_ ), .A2(\mreg/_04569_ ), .A3(\mreg/_02447_ ), .ZN(\mreg/_03537_ ) );
NAND2_X1 \mreg/_09467_ ( .A1(\mreg/_03536_ ), .A2(\mreg/_03537_ ), .ZN(\mreg/_03538_ ) );
AOI221_X4 \mreg/_09468_ ( .A(\mreg/_03538_ ), .B1(\mreg/_02227_ ), .B2(\mreg/_02550_ ), .C1(\mreg/_04665_ ), .C2(\mreg/_02603_ ), .ZN(\mreg/_03539_ ) );
NAND4_X1 \mreg/_09469_ ( .A1(\mreg/_02585_ ), .A2(\mreg/_02644_ ), .A3(\mreg/_04505_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03540_ ) );
OAI21_X1 \mreg/_09470_ ( .A(\mreg/_03540_ ), .B1(\mreg/_02539_ ), .B2(\mreg/_02231_ ), .ZN(\mreg/_03541_ ) );
AOI221_X4 \mreg/_09471_ ( .A(\mreg/_03541_ ), .B1(\mreg/_04473_ ), .B2(\mreg/_02542_ ), .C1(\mreg/_04441_ ), .C2(\mreg/_02544_ ), .ZN(\mreg/_03542_ ) );
NAND3_X1 \mreg/_09472_ ( .A1(\mreg/_02845_ ), .A2(\mreg/_04185_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03543_ ) );
NAND3_X1 \mreg/_09473_ ( .A1(\mreg/_02511_ ), .A2(\mreg/_04153_ ), .A3(\mreg/_02581_ ), .ZN(\mreg/_03544_ ) );
NAND4_X1 \mreg/_09474_ ( .A1(\mreg/_02587_ ), .A2(\mreg/_04217_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02581_ ), .ZN(\mreg/_03545_ ) );
NAND4_X1 \mreg/_09475_ ( .A1(\mreg/_02589_ ), .A2(\mreg/_02581_ ), .A3(\mreg/_04249_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03546_ ) );
NAND4_X1 \mreg/_09476_ ( .A1(\mreg/_03543_ ), .A2(\mreg/_03544_ ), .A3(\mreg/_03545_ ), .A4(\mreg/_03546_ ), .ZN(\mreg/_03547_ ) );
NAND3_X1 \mreg/_09477_ ( .A1(\mreg/_02455_ ), .A2(\mreg/_04377_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03548_ ) );
NAND3_X1 \mreg/_09478_ ( .A1(\mreg/_02842_ ), .A2(\mreg/_04409_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03549_ ) );
NAND2_X1 \mreg/_09479_ ( .A1(\mreg/_03548_ ), .A2(\mreg/_03549_ ), .ZN(\mreg/_03550_ ) );
AND3_X1 \mreg/_09480_ ( .A1(\mreg/_02503_ ), .A2(\mreg/_04345_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03551_ ) );
AND3_X1 \mreg/_09481_ ( .A1(\mreg/_02837_ ), .A2(\mreg/_04313_ ), .A3(\mreg/_02512_ ), .ZN(\mreg/_03552_ ) );
NOR4_X1 \mreg/_09482_ ( .A1(\mreg/_03547_ ), .A2(\mreg/_03550_ ), .A3(\mreg/_03551_ ), .A4(\mreg/_03552_ ), .ZN(\mreg/_03553_ ) );
NAND4_X1 \mreg/_09483_ ( .A1(\mreg/_03535_ ), .A2(\mreg/_03539_ ), .A3(\mreg/_03542_ ), .A4(\mreg/_03553_ ), .ZN(\mreg/_03897_ ) );
NAND3_X1 \mreg/_09484_ ( .A1(\mreg/_02531_ ), .A2(\mreg/_04570_ ), .A3(\mreg/_02533_ ), .ZN(\mreg/_03554_ ) );
NAND4_X1 \mreg/_09485_ ( .A1(\mreg/_03015_ ), .A2(\mreg/_02879_ ), .A3(\mreg/_04506_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03555_ ) );
OAI21_X1 \mreg/_09486_ ( .A(\mreg/_03555_ ), .B1(\mreg/_02538_ ), .B2(\mreg/_02268_ ), .ZN(\mreg/_03556_ ) );
AOI221_X4 \mreg/_09487_ ( .A(\mreg/_03556_ ), .B1(\mreg/_04474_ ), .B2(\mreg/_02541_ ), .C1(\mreg/_04442_ ), .C2(\mreg/_02543_ ), .ZN(\mreg/_03557_ ) );
NAND3_X1 \mreg/_09488_ ( .A1(\mreg/_02546_ ), .A2(\mreg/_04602_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03558_ ) );
AND3_X1 \mreg/_09489_ ( .A1(\mreg/_02571_ ), .A2(\mreg/_04666_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03559_ ) );
AOI21_X1 \mreg/_09490_ ( .A(\mreg/_03559_ ), .B1(\mreg/_02264_ ), .B2(\mreg/_02550_ ), .ZN(\mreg/_03560_ ) );
AND4_X1 \mreg/_09491_ ( .A1(\mreg/_03554_ ), .A2(\mreg/_03557_ ), .A3(\mreg/_03558_ ), .A4(\mreg/_03560_ ), .ZN(\mreg/_03561_ ) );
NAND3_X1 \mreg/_09492_ ( .A1(\mreg/_02672_ ), .A2(\mreg/_04378_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03562_ ) );
NAND4_X1 \mreg/_09493_ ( .A1(\mreg/_02451_ ), .A2(\mreg/_04218_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02499_ ), .ZN(\mreg/_03563_ ) );
OAI21_X1 \mreg/_09494_ ( .A(\mreg/_03563_ ), .B1(\mreg/_02492_ ), .B2(\mreg/_02276_ ), .ZN(\mreg/_03564_ ) );
AOI221_X4 \mreg/_09495_ ( .A(\mreg/_03564_ ), .B1(\mreg/_04186_ ), .B2(\mreg/_02495_ ), .C1(\mreg/_04154_ ), .C2(\mreg/_02500_ ), .ZN(\mreg/_03565_ ) );
NAND3_X1 \mreg/_09496_ ( .A1(\mreg/_02508_ ), .A2(\mreg/_04410_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03566_ ) );
AND3_X1 \mreg/_09497_ ( .A1(\mreg/_02520_ ), .A2(\mreg/_04314_ ), .A3(\mreg/_02466_ ), .ZN(\mreg/_03567_ ) );
AOI21_X1 \mreg/_09498_ ( .A(\mreg/_03567_ ), .B1(\mreg/_04346_ ), .B2(\mreg/_02947_ ), .ZN(\mreg/_03568_ ) );
AND4_X1 \mreg/_09499_ ( .A1(\mreg/_03562_ ), .A2(\mreg/_03565_ ), .A3(\mreg/_03566_ ), .A4(\mreg/_03568_ ), .ZN(\mreg/_03569_ ) );
NAND3_X1 \mreg/_09500_ ( .A1(\mreg/_02583_ ), .A2(\mreg/_04282_ ), .A3(\mreg/_02820_ ), .ZN(\mreg/_03570_ ) );
AND3_X1 \mreg/_09501_ ( .A1(\mreg/_02632_ ), .A2(\mreg/_04858_ ), .A3(\mreg/_02572_ ), .ZN(\mreg/_03571_ ) );
AOI21_X1 \mreg/_09502_ ( .A(\mreg/_03571_ ), .B1(\mreg/_04826_ ), .B2(\mreg/_02636_ ), .ZN(\mreg/_03572_ ) );
AOI22_X1 \mreg/_09503_ ( .A1(\mreg/_04634_ ), .A2(\mreg/_02724_ ), .B1(\mreg/_02723_ ), .B2(\mreg/_04730_ ), .ZN(\mreg/_03573_ ) );
AOI22_X1 \mreg/_09504_ ( .A1(\mreg/_02814_ ), .A2(\mreg/_04794_ ), .B1(\mreg/_04762_ ), .B2(\mreg/_02817_ ), .ZN(\mreg/_03574_ ) );
AND4_X1 \mreg/_09505_ ( .A1(\mreg/_03570_ ), .A2(\mreg/_03572_ ), .A3(\mreg/_03573_ ), .A4(\mreg/_03574_ ), .ZN(\mreg/_03575_ ) );
NAND3_X1 \mreg/_09506_ ( .A1(\mreg/_02641_ ), .A2(\mreg/_03962_ ), .A3(\mreg/_02642_ ), .ZN(\mreg/_03576_ ) );
NAND3_X1 \mreg/_09507_ ( .A1(\mreg/_02445_ ), .A2(\mreg/_04026_ ), .A3(\mreg/_02448_ ), .ZN(\mreg/_03577_ ) );
NAND3_X1 \mreg/_09508_ ( .A1(\mreg/_02571_ ), .A2(\mreg/_04090_ ), .A3(\mreg/_02566_ ), .ZN(\mreg/_03578_ ) );
NAND3_X1 \mreg/_09509_ ( .A1(\mreg/_02696_ ), .A2(\mreg/_04058_ ), .A3(\mreg/_02572_ ), .ZN(\mreg/_03579_ ) );
NAND3_X1 \mreg/_09510_ ( .A1(\mreg/_02699_ ), .A2(\mreg/_04122_ ), .A3(\mreg/_02633_ ), .ZN(\mreg/_03580_ ) );
AND4_X1 \mreg/_09511_ ( .A1(\mreg/_03577_ ), .A2(\mreg/_03578_ ), .A3(\mreg/_03579_ ), .A4(\mreg/_03580_ ), .ZN(\mreg/_03581_ ) );
NAND3_X1 \mreg/_09512_ ( .A1(\mreg/_02647_ ), .A2(\mreg/_03994_ ), .A3(\mreg/_02648_ ), .ZN(\mreg/_03582_ ) );
NAND3_X1 \mreg/_09513_ ( .A1(\mreg/_02472_ ), .A2(\mreg/_04922_ ), .A3(\mreg/_02428_ ), .ZN(\mreg/_03583_ ) );
NAND3_X1 \mreg/_09514_ ( .A1(\mreg/_02629_ ), .A2(\mreg/_02851_ ), .A3(\mreg/_04890_ ), .ZN(\mreg/_03584_ ) );
AND2_X1 \mreg/_09515_ ( .A1(\mreg/_03583_ ), .A2(\mreg/_03584_ ), .ZN(\mreg/_03585_ ) );
AND4_X1 \mreg/_09516_ ( .A1(\mreg/_03576_ ), .A2(\mreg/_03581_ ), .A3(\mreg/_03582_ ), .A4(\mreg/_03585_ ), .ZN(\mreg/_03586_ ) );
NAND4_X1 \mreg/_09517_ ( .A1(\mreg/_03561_ ), .A2(\mreg/_03569_ ), .A3(\mreg/_03575_ ), .A4(\mreg/_03586_ ), .ZN(\mreg/_03898_ ) );
NAND3_X1 \mreg/_09518_ ( .A1(\mreg/_02672_ ), .A2(\mreg/_04379_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03587_ ) );
NAND4_X1 \mreg/_09519_ ( .A1(\mreg/_03015_ ), .A2(\mreg/_04219_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02609_ ), .ZN(\mreg/_03588_ ) );
OAI21_X1 \mreg/_09520_ ( .A(\mreg/_03588_ ), .B1(\mreg/_02611_ ), .B2(\mreg/_02310_ ), .ZN(\mreg/_03589_ ) );
AOI221_X4 \mreg/_09521_ ( .A(\mreg/_03589_ ), .B1(\mreg/_04187_ ), .B2(\mreg/_02496_ ), .C1(\mreg/_04155_ ), .C2(\mreg/_02614_ ), .ZN(\mreg/_03590_ ) );
NAND3_X1 \mreg/_09522_ ( .A1(\mreg/_02674_ ), .A2(\mreg/_04411_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03591_ ) );
AND3_X1 \mreg/_09523_ ( .A1(\mreg/_02767_ ), .A2(\mreg/_04347_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03592_ ) );
AOI21_X1 \mreg/_09524_ ( .A(\mreg/_03592_ ), .B1(\mreg/_04315_ ), .B2(\mreg/_02807_ ), .ZN(\mreg/_03593_ ) );
AND4_X1 \mreg/_09525_ ( .A1(\mreg/_03587_ ), .A2(\mreg/_03590_ ), .A3(\mreg/_03591_ ), .A4(\mreg/_03593_ ), .ZN(\mreg/_03594_ ) );
NAND3_X1 \mreg/_09526_ ( .A1(\mreg/_02531_ ), .A2(\mreg/_04571_ ), .A3(\mreg/_02533_ ), .ZN(\mreg/_03595_ ) );
NAND3_X1 \mreg/_09527_ ( .A1(\mreg/_02516_ ), .A2(\mreg/_04667_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03596_ ) );
NAND3_X1 \mreg/_09528_ ( .A1(\mreg/_02546_ ), .A2(\mreg/_04603_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03597_ ) );
NAND3_X1 \mreg/_09529_ ( .A1(\mreg/_02524_ ), .A2(\mreg/_02299_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03598_ ) );
AND4_X1 \mreg/_09530_ ( .A1(\mreg/_03595_ ), .A2(\mreg/_03596_ ), .A3(\mreg/_03597_ ), .A4(\mreg/_03598_ ), .ZN(\mreg/_03599_ ) );
AND4_X1 \mreg/_09531_ ( .A1(\mreg/_04507_ ), .A2(\mreg/_02585_ ), .A3(\mreg/_02536_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03600_ ) );
AND4_X1 \mreg/_09532_ ( .A1(\mreg/_04539_ ), .A2(\mreg/_02536_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02413_ ), .ZN(\mreg/_03601_ ) );
OR2_X1 \mreg/_09533_ ( .A1(\mreg/_03600_ ), .A2(\mreg/_03601_ ), .ZN(\mreg/_03602_ ) );
AOI221_X4 \mreg/_09534_ ( .A(\mreg/_03602_ ), .B1(\mreg/_04475_ ), .B2(\mreg/_02542_ ), .C1(\mreg/_04443_ ), .C2(\mreg/_02544_ ), .ZN(\mreg/_03603_ ) );
AND3_X1 \mreg/_09535_ ( .A1(\mreg/_02855_ ), .A2(\mreg/_04731_ ), .A3(\mreg/_02415_ ), .ZN(\mreg/_03604_ ) );
AOI221_X4 \mreg/_09536_ ( .A(\mreg/_03604_ ), .B1(\mreg/_02627_ ), .B2(\mreg/_04635_ ), .C1(\mreg/_04283_ ), .C2(\mreg/_02420_ ), .ZN(\mreg/_03605_ ) );
NAND3_X1 \mreg/_09537_ ( .A1(\mreg/_02463_ ), .A2(\mreg/_04795_ ), .A3(\mreg/_02460_ ), .ZN(\mreg/_03606_ ) );
NAND3_X1 \mreg/_09538_ ( .A1(\mreg/_02454_ ), .A2(\mreg/_04827_ ), .A3(\mreg/_02566_ ), .ZN(\mreg/_03607_ ) );
NAND3_X1 \mreg/_09539_ ( .A1(\mreg/_02632_ ), .A2(\mreg/_04859_ ), .A3(\mreg/_02688_ ), .ZN(\mreg/_03608_ ) );
NAND3_X1 \mreg/_09540_ ( .A1(\mreg/_02684_ ), .A2(\mreg/_02568_ ), .A3(\mreg/_04763_ ), .ZN(\mreg/_03609_ ) );
AND4_X1 \mreg/_09541_ ( .A1(\mreg/_03606_ ), .A2(\mreg/_03607_ ), .A3(\mreg/_03608_ ), .A4(\mreg/_03609_ ), .ZN(\mreg/_03610_ ) );
NAND3_X1 \mreg/_09542_ ( .A1(\mreg/_02471_ ), .A2(\mreg/_04923_ ), .A3(\mreg/_02464_ ), .ZN(\mreg/_03611_ ) );
NAND3_X1 \mreg/_09543_ ( .A1(\mreg/_02476_ ), .A2(\mreg/_03963_ ), .A3(\mreg/_02688_ ), .ZN(\mreg/_03612_ ) );
NAND3_X1 \mreg/_09544_ ( .A1(\mreg/_02729_ ), .A2(\mreg/_02644_ ), .A3(\mreg/_04891_ ), .ZN(\mreg/_03613_ ) );
NAND3_X1 \mreg/_09545_ ( .A1(\mreg/_02484_ ), .A2(\mreg/_03995_ ), .A3(\mreg/_02697_ ), .ZN(\mreg/_03614_ ) );
AND4_X1 \mreg/_09546_ ( .A1(\mreg/_03611_ ), .A2(\mreg/_03612_ ), .A3(\mreg/_03613_ ), .A4(\mreg/_03614_ ), .ZN(\mreg/_03615_ ) );
NAND3_X1 \mreg/_09547_ ( .A1(\mreg/_02479_ ), .A2(\mreg/_04027_ ), .A3(\mreg/_02447_ ), .ZN(\mreg/_03616_ ) );
NAND3_X1 \mreg/_09548_ ( .A1(\mreg/_02431_ ), .A2(\mreg/_04091_ ), .A3(\mreg/_02691_ ), .ZN(\mreg/_03617_ ) );
NAND3_X1 \mreg/_09549_ ( .A1(\mreg/_02440_ ), .A2(\mreg/_04059_ ), .A3(\mreg/_02697_ ), .ZN(\mreg/_03618_ ) );
NAND3_X1 \mreg/_09550_ ( .A1(\mreg/_02425_ ), .A2(\mreg/_04123_ ), .A3(\mreg/_02700_ ), .ZN(\mreg/_03619_ ) );
AND4_X1 \mreg/_09551_ ( .A1(\mreg/_03616_ ), .A2(\mreg/_03617_ ), .A3(\mreg/_03618_ ), .A4(\mreg/_03619_ ), .ZN(\mreg/_03620_ ) );
AND4_X2 \mreg/_09552_ ( .A1(\mreg/_03605_ ), .A2(\mreg/_03610_ ), .A3(\mreg/_03615_ ), .A4(\mreg/_03620_ ), .ZN(\mreg/_03621_ ) );
NAND4_X1 \mreg/_09553_ ( .A1(\mreg/_03594_ ), .A2(\mreg/_03599_ ), .A3(\mreg/_03603_ ), .A4(\mreg/_03621_ ), .ZN(\mreg/_03899_ ) );
AOI22_X1 \mreg/_09554_ ( .A1(\mreg/_04829_ ), .A2(\mreg/_02635_ ), .B1(\mreg/_02814_ ), .B2(\mreg/_04797_ ), .ZN(\mreg/_03622_ ) );
NAND3_X1 \mreg/_09555_ ( .A1(\mreg/_02741_ ), .A2(\mreg/_02512_ ), .A3(\mreg/_04765_ ), .ZN(\mreg/_03623_ ) );
OAI211_X2 \mreg/_09556_ ( .A(\mreg/_03622_ ), .B(\mreg/_03623_ ), .C1(\mreg/_02359_ ), .C2(\mreg/_03112_ ), .ZN(\mreg/_03624_ ) );
AND3_X1 \mreg/_09557_ ( .A1(\mreg/_02431_ ), .A2(\mreg/_04669_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03625_ ) );
AND3_X1 \mreg/_09558_ ( .A1(\mreg/_02462_ ), .A2(\mreg/_04349_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03626_ ) );
AND3_X4 \mreg/_09559_ ( .A1(\mreg/_02498_ ), .A2(\mreg/_04317_ ), .A3(\mreg/_02452_ ), .ZN(\mreg/_03627_ ) );
AND4_X1 \mreg/_09560_ ( .A1(\mreg/_04221_ ), .A2(\mreg/_02451_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02407_ ), .ZN(\mreg/_03628_ ) );
AND4_X4 \mreg/_09561_ ( .A1(\mreg/_04253_ ), .A2(\mreg/_02413_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02407_ ), .ZN(\mreg/_03629_ ) );
OR4_X4 \mreg/_09562_ ( .A1(\mreg/_03626_ ), .A2(\mreg/_03627_ ), .A3(\mreg/_03628_ ), .A4(\mreg/_03629_ ), .ZN(\mreg/_03630_ ) );
AND3_X1 \mreg/_09563_ ( .A1(\mreg/_02425_ ), .A2(\mreg/_02335_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03631_ ) );
NAND4_X1 \mreg/_09564_ ( .A1(\mreg/_02585_ ), .A2(\mreg/_02480_ ), .A3(\mreg/_04509_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03632_ ) );
OAI21_X1 \mreg/_09565_ ( .A(\mreg/_03632_ ), .B1(\mreg/_02539_ ), .B2(\mreg/_02362_ ), .ZN(\mreg/_03633_ ) );
OR4_X4 \mreg/_09566_ ( .A1(\mreg/_03625_ ), .A2(\mreg/_03630_ ), .A3(\mreg/_03631_ ), .A4(\mreg/_03633_ ), .ZN(\mreg/_03634_ ) );
AOI22_X1 \mreg/_09567_ ( .A1(\mreg/_02560_ ), .A2(\mreg/_03965_ ), .B1(\mreg/_02734_ ), .B2(\mreg/_04925_ ), .ZN(\mreg/_03635_ ) );
NAND3_X1 \mreg/_09568_ ( .A1(\mreg/_02426_ ), .A2(\mreg/_04125_ ), .A3(\mreg/_02623_ ), .ZN(\mreg/_03636_ ) );
OAI211_X2 \mreg/_09569_ ( .A(\mreg/_03635_ ), .B(\mreg/_03636_ ), .C1(\mreg/_02368_ ), .C2(\mreg/_03116_ ), .ZN(\mreg/_03637_ ) );
NAND3_X1 \mreg/_09570_ ( .A1(\mreg/_02458_ ), .A2(\mreg/_04861_ ), .A3(\mreg/_02433_ ), .ZN(\mreg/_03638_ ) );
NAND3_X1 \mreg/_09571_ ( .A1(\mreg/_02419_ ), .A2(\mreg/_04285_ ), .A3(\mreg/_02433_ ), .ZN(\mreg/_03639_ ) );
NAND3_X1 \mreg/_09572_ ( .A1(\mreg/_02409_ ), .A2(\mreg/_04637_ ), .A3(\mreg/_02433_ ), .ZN(\mreg/_03640_ ) );
NAND3_X1 \mreg/_09573_ ( .A1(\mreg/_02444_ ), .A2(\mreg/_02480_ ), .A3(\mreg/_04893_ ), .ZN(\mreg/_03641_ ) );
NAND4_X1 \mreg/_09574_ ( .A1(\mreg/_03638_ ), .A2(\mreg/_03639_ ), .A3(\mreg/_03640_ ), .A4(\mreg/_03641_ ), .ZN(\mreg/_03642_ ) );
NAND3_X1 \mreg/_09575_ ( .A1(\mreg/_02443_ ), .A2(\mreg/_04029_ ), .A3(\mreg/_02446_ ), .ZN(\mreg/_03643_ ) );
OAI221_X1 \mreg/_09576_ ( .A(\mreg/_03643_ ), .B1(\mreg/_02749_ ), .B2(\mreg/_02347_ ), .C1(\mreg/_02348_ ), .C2(\mreg/_02739_ ), .ZN(\mreg/_03644_ ) );
NAND3_X1 \mreg/_09577_ ( .A1(\mreg/_02470_ ), .A2(\mreg/_04477_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03645_ ) );
NAND3_X1 \mreg/_09578_ ( .A1(\mreg/_02597_ ), .A2(\mreg/_04605_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03646_ ) );
NAND3_X1 \mreg/_09579_ ( .A1(\mreg/_02599_ ), .A2(\mreg/_04573_ ), .A3(\mreg/_02446_ ), .ZN(\mreg/_03647_ ) );
NAND3_X1 \mreg/_09580_ ( .A1(\mreg/_02599_ ), .A2(\mreg/_04445_ ), .A3(\mreg/_02536_ ), .ZN(\mreg/_03648_ ) );
NAND4_X1 \mreg/_09581_ ( .A1(\mreg/_03645_ ), .A2(\mreg/_03646_ ), .A3(\mreg/_03647_ ), .A4(\mreg/_03648_ ), .ZN(\mreg/_03649_ ) );
NAND3_X1 \mreg/_09582_ ( .A1(\mreg/_02453_ ), .A2(\mreg/_04381_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03650_ ) );
NAND3_X4 \mreg/_09583_ ( .A1(\mreg/_02458_ ), .A2(\mreg/_04413_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03651_ ) );
NAND3_X1 \mreg/_09584_ ( .A1(\mreg/_02599_ ), .A2(\mreg/_04157_ ), .A3(\mreg/_02579_ ), .ZN(\mreg/_03652_ ) );
NAND3_X1 \mreg/_09585_ ( .A1(\mreg/_02419_ ), .A2(\mreg/_04189_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03653_ ) );
NAND4_X1 \mreg/_09586_ ( .A1(\mreg/_03650_ ), .A2(\mreg/_03651_ ), .A3(\mreg/_03652_ ), .A4(\mreg/_03653_ ), .ZN(\mreg/_03654_ ) );
OR4_X2 \mreg/_09587_ ( .A1(\mreg/_03642_ ), .A2(\mreg/_03644_ ), .A3(\mreg/_03649_ ), .A4(\mreg/_03654_ ), .ZN(\mreg/_03655_ ) );
OR4_X2 \mreg/_09588_ ( .A1(\mreg/_03624_ ), .A2(\mreg/_03634_ ), .A3(\mreg/_03637_ ), .A4(\mreg/_03655_ ), .ZN(\mreg/_03901_ ) );
NAND3_X1 \mreg/_09589_ ( .A1(\mreg/_02516_ ), .A2(\mreg/_04670_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03656_ ) );
NAND4_X1 \mreg/_09590_ ( .A1(\mreg/_02608_ ), .A2(\mreg/_02474_ ), .A3(\mreg/_04510_ ), .A4(\mreg/_03872_ ), .ZN(\mreg/_03657_ ) );
OAI21_X1 \mreg/_09591_ ( .A(\mreg/_03657_ ), .B1(\mreg/_02538_ ), .B2(\mreg/_02377_ ), .ZN(\mreg/_03658_ ) );
AOI221_X4 \mreg/_09592_ ( .A(\mreg/_03658_ ), .B1(\mreg/_04478_ ), .B2(\mreg/_02541_ ), .C1(\mreg/_04446_ ), .C2(\mreg/_02543_ ), .ZN(\mreg/_03659_ ) );
NAND3_X1 \mreg/_09593_ ( .A1(\mreg/_02524_ ), .A2(\mreg/_02374_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03660_ ) );
AND3_X1 \mreg/_09594_ ( .A1(\mreg/_02619_ ), .A2(\mreg/_04574_ ), .A3(\mreg/_02664_ ), .ZN(\mreg/_03661_ ) );
AOI21_X1 \mreg/_09595_ ( .A(\mreg/_03661_ ), .B1(\mreg/_02527_ ), .B2(\mreg/_04606_ ), .ZN(\mreg/_03662_ ) );
AND4_X1 \mreg/_09596_ ( .A1(\mreg/_03656_ ), .A2(\mreg/_03659_ ), .A3(\mreg/_03660_ ), .A4(\mreg/_03662_ ), .ZN(\mreg/_03663_ ) );
NAND4_X1 \mreg/_09597_ ( .A1(\mreg/_02586_ ), .A2(\mreg/_04222_ ), .A3(\mreg/_03872_ ), .A4(\mreg/_02579_ ), .ZN(\mreg/_03664_ ) );
OAI21_X1 \mreg/_09598_ ( .A(\mreg/_03664_ ), .B1(\mreg/_02493_ ), .B2(\mreg/_02385_ ), .ZN(\mreg/_03665_ ) );
AOI221_X4 \mreg/_09599_ ( .A(\mreg/_03665_ ), .B1(\mreg/_04190_ ), .B2(\mreg/_02496_ ), .C1(\mreg/_04158_ ), .C2(\mreg/_02501_ ), .ZN(\mreg/_03666_ ) );
NAND3_X1 \mreg/_09600_ ( .A1(\mreg/_02506_ ), .A2(\mreg/_04382_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03667_ ) );
NAND3_X1 \mreg/_09601_ ( .A1(\mreg/_02674_ ), .A2(\mreg/_04414_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03668_ ) );
NAND3_X1 \mreg/_09602_ ( .A1(\mreg/_02504_ ), .A2(\mreg/_04350_ ), .A3(\mreg/_03872_ ), .ZN(\mreg/_03669_ ) );
NAND3_X1 \mreg/_09603_ ( .A1(\mreg/_02511_ ), .A2(\mreg/_04318_ ), .A3(\mreg/_02513_ ), .ZN(\mreg/_03670_ ) );
AND4_X1 \mreg/_09604_ ( .A1(\mreg/_03667_ ), .A2(\mreg/_03668_ ), .A3(\mreg/_03669_ ), .A4(\mreg/_03670_ ), .ZN(\mreg/_03671_ ) );
AND3_X1 \mreg/_09605_ ( .A1(\mreg/_02414_ ), .A2(\mreg/_04734_ ), .A3(\mreg/_02415_ ), .ZN(\mreg/_03672_ ) );
AOI221_X4 \mreg/_09606_ ( .A(\mreg/_03672_ ), .B1(\mreg/_02627_ ), .B2(\mreg/_04638_ ), .C1(\mreg/_04286_ ), .C2(\mreg/_02420_ ), .ZN(\mreg/_03673_ ) );
NAND3_X1 \mreg/_09607_ ( .A1(\mreg/_02463_ ), .A2(\mreg/_04798_ ), .A3(\mreg/_02460_ ), .ZN(\mreg/_03674_ ) );
NAND3_X1 \mreg/_09608_ ( .A1(\mreg/_02454_ ), .A2(\mreg/_04830_ ), .A3(\mreg/_02566_ ), .ZN(\mreg/_03675_ ) );
NAND3_X1 \mreg/_09609_ ( .A1(\mreg/_02632_ ), .A2(\mreg/_04862_ ), .A3(\mreg/_02688_ ), .ZN(\mreg/_03676_ ) );
NAND3_X1 \mreg/_09610_ ( .A1(\mreg/_02684_ ), .A2(\mreg/_02568_ ), .A3(\mreg/_04766_ ), .ZN(\mreg/_03677_ ) );
AND4_X1 \mreg/_09611_ ( .A1(\mreg/_03674_ ), .A2(\mreg/_03675_ ), .A3(\mreg/_03676_ ), .A4(\mreg/_03677_ ), .ZN(\mreg/_03678_ ) );
NAND3_X1 \mreg/_09612_ ( .A1(\mreg/_02471_ ), .A2(\mreg/_04926_ ), .A3(\mreg/_02563_ ), .ZN(\mreg/_03679_ ) );
NAND3_X1 \mreg/_09613_ ( .A1(\mreg/_02476_ ), .A2(\mreg/_03966_ ), .A3(\mreg/_02688_ ), .ZN(\mreg/_03680_ ) );
NAND3_X1 \mreg/_09614_ ( .A1(\mreg/_02729_ ), .A2(\mreg/_02644_ ), .A3(\mreg/_04894_ ), .ZN(\mreg/_03681_ ) );
NAND3_X1 \mreg/_09615_ ( .A1(\mreg/_02484_ ), .A2(\mreg/_03998_ ), .A3(\mreg/_02697_ ), .ZN(\mreg/_03682_ ) );
AND4_X1 \mreg/_09616_ ( .A1(\mreg/_03679_ ), .A2(\mreg/_03680_ ), .A3(\mreg/_03681_ ), .A4(\mreg/_03682_ ), .ZN(\mreg/_03683_ ) );
NAND3_X1 \mreg/_09617_ ( .A1(\mreg/_02479_ ), .A2(\mreg/_04030_ ), .A3(\mreg/_02447_ ), .ZN(\mreg/_03684_ ) );
NAND3_X1 \mreg/_09618_ ( .A1(\mreg/_02431_ ), .A2(\mreg/_04094_ ), .A3(\mreg/_02691_ ), .ZN(\mreg/_03685_ ) );
NAND3_X1 \mreg/_09619_ ( .A1(\mreg/_02440_ ), .A2(\mreg/_04062_ ), .A3(\mreg/_02697_ ), .ZN(\mreg/_03686_ ) );
NAND3_X1 \mreg/_09620_ ( .A1(\mreg/_02425_ ), .A2(\mreg/_04126_ ), .A3(\mreg/_02700_ ), .ZN(\mreg/_03687_ ) );
AND4_X1 \mreg/_09621_ ( .A1(\mreg/_03684_ ), .A2(\mreg/_03685_ ), .A3(\mreg/_03686_ ), .A4(\mreg/_03687_ ), .ZN(\mreg/_03688_ ) );
AND4_X1 \mreg/_09622_ ( .A1(\mreg/_03673_ ), .A2(\mreg/_03678_ ), .A3(\mreg/_03683_ ), .A4(\mreg/_03688_ ), .ZN(\mreg/_03689_ ) );
NAND4_X1 \mreg/_09623_ ( .A1(\mreg/_03663_ ), .A2(\mreg/_03666_ ), .A3(\mreg/_03671_ ), .A4(\mreg/_03689_ ), .ZN(\mreg/_03902_ ) );
NOR2_X4 \mreg/_09624_ ( .A1(\mreg/_04936_ ), .A2(\mreg/_04937_ ), .ZN(\mreg/_03690_ ) );
NOR2_X4 \mreg/_09625_ ( .A1(\mreg/_04934_ ), .A2(\mreg/_04935_ ), .ZN(\mreg/_03691_ ) );
INV_X1 \mreg/_09626_ ( .A(\mreg/_04938_ ), .ZN(\mreg/_03692_ ) );
NAND3_X1 \mreg/_09627_ ( .A1(\mreg/_03690_ ), .A2(\mreg/_03691_ ), .A3(\mreg/_03692_ ), .ZN(\mreg/_03693_ ) );
AND2_X1 \mreg/_09628_ ( .A1(\mreg/_04971_ ), .A2(\mreg/_01054_ ), .ZN(\mreg/_03694_ ) );
NAND2_X1 \mreg/_09629_ ( .A1(\mreg/_03693_ ), .A2(\mreg/_03694_ ), .ZN(\mreg/_03695_ ) );
BUF_X4 \mreg/_09630_ ( .A(\mreg/_03695_ ), .Z(\mreg/_03696_ ) );
NAND2_X1 \mreg/_09631_ ( .A1(\mreg/_04936_ ), .A2(\mreg/_04937_ ), .ZN(\mreg/_03697_ ) );
NAND2_X1 \mreg/_09632_ ( .A1(\mreg/_04934_ ), .A2(\mreg/_04935_ ), .ZN(\mreg/_03698_ ) );
NOR2_X1 \mreg/_09633_ ( .A1(\mreg/_03697_ ), .A2(\mreg/_03698_ ), .ZN(\mreg/_03699_ ) );
NAND2_X1 \mreg/_09634_ ( .A1(\mreg/_03699_ ), .A2(\mreg/_04938_ ), .ZN(\mreg/_03700_ ) );
NOR2_X1 \mreg/_09635_ ( .A1(\mreg/_03696_ ), .A2(\mreg/_03700_ ), .ZN(\mreg/_03701_ ) );
BUF_X4 \mreg/_09636_ ( .A(\mreg/_03701_ ), .Z(\mreg/_03702_ ) );
MUX2_X1 \mreg/_09637_ ( .A(\mreg/_04678_ ), .B(\mreg/_04939_ ), .S(\mreg/_03702_ ), .Z(\mreg/_00062_ ) );
MUX2_X1 \mreg/_09638_ ( .A(\mreg/_04689_ ), .B(\mreg/_04950_ ), .S(\mreg/_03702_ ), .Z(\mreg/_00063_ ) );
MUX2_X1 \mreg/_09639_ ( .A(\mreg/_04700_ ), .B(\mreg/_04961_ ), .S(\mreg/_03702_ ), .Z(\mreg/_00064_ ) );
MUX2_X1 \mreg/_09640_ ( .A(\mreg/_04703_ ), .B(\mreg/_04964_ ), .S(\mreg/_03702_ ), .Z(\mreg/_00065_ ) );
MUX2_X1 \mreg/_09641_ ( .A(\mreg/_04704_ ), .B(\mreg/_04965_ ), .S(\mreg/_03702_ ), .Z(\mreg/_00066_ ) );
MUX2_X1 \mreg/_09642_ ( .A(\mreg/_04705_ ), .B(\mreg/_04966_ ), .S(\mreg/_03702_ ), .Z(\mreg/_00067_ ) );
MUX2_X1 \mreg/_09643_ ( .A(\mreg/_04706_ ), .B(\mreg/_04967_ ), .S(\mreg/_03702_ ), .Z(\mreg/_00068_ ) );
MUX2_X1 \mreg/_09644_ ( .A(\mreg/_04707_ ), .B(\mreg/_04968_ ), .S(\mreg/_03702_ ), .Z(\mreg/_00069_ ) );
MUX2_X1 \mreg/_09645_ ( .A(\mreg/_04708_ ), .B(\mreg/_04969_ ), .S(\mreg/_03702_ ), .Z(\mreg/_00070_ ) );
MUX2_X1 \mreg/_09646_ ( .A(\mreg/_04709_ ), .B(\mreg/_04970_ ), .S(\mreg/_03702_ ), .Z(\mreg/_00071_ ) );
BUF_X4 \mreg/_09647_ ( .A(\mreg/_03701_ ), .Z(\mreg/_03703_ ) );
MUX2_X1 \mreg/_09648_ ( .A(\mreg/_04679_ ), .B(\mreg/_04940_ ), .S(\mreg/_03703_ ), .Z(\mreg/_00072_ ) );
MUX2_X1 \mreg/_09649_ ( .A(\mreg/_04680_ ), .B(\mreg/_04941_ ), .S(\mreg/_03703_ ), .Z(\mreg/_00073_ ) );
MUX2_X1 \mreg/_09650_ ( .A(\mreg/_04681_ ), .B(\mreg/_04942_ ), .S(\mreg/_03703_ ), .Z(\mreg/_00074_ ) );
MUX2_X1 \mreg/_09651_ ( .A(\mreg/_04682_ ), .B(\mreg/_04943_ ), .S(\mreg/_03703_ ), .Z(\mreg/_00075_ ) );
MUX2_X1 \mreg/_09652_ ( .A(\mreg/_04683_ ), .B(\mreg/_04944_ ), .S(\mreg/_03703_ ), .Z(\mreg/_00076_ ) );
MUX2_X1 \mreg/_09653_ ( .A(\mreg/_04684_ ), .B(\mreg/_04945_ ), .S(\mreg/_03703_ ), .Z(\mreg/_00077_ ) );
MUX2_X1 \mreg/_09654_ ( .A(\mreg/_04685_ ), .B(\mreg/_04946_ ), .S(\mreg/_03703_ ), .Z(\mreg/_00078_ ) );
MUX2_X1 \mreg/_09655_ ( .A(\mreg/_04686_ ), .B(\mreg/_04947_ ), .S(\mreg/_03703_ ), .Z(\mreg/_00079_ ) );
MUX2_X1 \mreg/_09656_ ( .A(\mreg/_04687_ ), .B(\mreg/_04948_ ), .S(\mreg/_03703_ ), .Z(\mreg/_00080_ ) );
MUX2_X1 \mreg/_09657_ ( .A(\mreg/_04688_ ), .B(\mreg/_04949_ ), .S(\mreg/_03703_ ), .Z(\mreg/_00081_ ) );
BUF_X4 \mreg/_09658_ ( .A(\mreg/_03701_ ), .Z(\mreg/_03704_ ) );
MUX2_X1 \mreg/_09659_ ( .A(\mreg/_04690_ ), .B(\mreg/_04951_ ), .S(\mreg/_03704_ ), .Z(\mreg/_00082_ ) );
MUX2_X1 \mreg/_09660_ ( .A(\mreg/_04691_ ), .B(\mreg/_04952_ ), .S(\mreg/_03704_ ), .Z(\mreg/_00083_ ) );
MUX2_X1 \mreg/_09661_ ( .A(\mreg/_04692_ ), .B(\mreg/_04953_ ), .S(\mreg/_03704_ ), .Z(\mreg/_00084_ ) );
MUX2_X1 \mreg/_09662_ ( .A(\mreg/_04693_ ), .B(\mreg/_04954_ ), .S(\mreg/_03704_ ), .Z(\mreg/_00085_ ) );
MUX2_X1 \mreg/_09663_ ( .A(\mreg/_04694_ ), .B(\mreg/_04955_ ), .S(\mreg/_03704_ ), .Z(\mreg/_00086_ ) );
MUX2_X1 \mreg/_09664_ ( .A(\mreg/_04695_ ), .B(\mreg/_04956_ ), .S(\mreg/_03704_ ), .Z(\mreg/_00087_ ) );
MUX2_X1 \mreg/_09665_ ( .A(\mreg/_04696_ ), .B(\mreg/_04957_ ), .S(\mreg/_03704_ ), .Z(\mreg/_00088_ ) );
MUX2_X1 \mreg/_09666_ ( .A(\mreg/_04697_ ), .B(\mreg/_04958_ ), .S(\mreg/_03704_ ), .Z(\mreg/_00089_ ) );
MUX2_X1 \mreg/_09667_ ( .A(\mreg/_04698_ ), .B(\mreg/_04959_ ), .S(\mreg/_03704_ ), .Z(\mreg/_00090_ ) );
MUX2_X1 \mreg/_09668_ ( .A(\mreg/_04699_ ), .B(\mreg/_04960_ ), .S(\mreg/_03704_ ), .Z(\mreg/_00091_ ) );
MUX2_X1 \mreg/_09669_ ( .A(\mreg/_04701_ ), .B(\mreg/_04962_ ), .S(\mreg/_03701_ ), .Z(\mreg/_00092_ ) );
MUX2_X1 \mreg/_09670_ ( .A(\mreg/_04702_ ), .B(\mreg/_04963_ ), .S(\mreg/_03701_ ), .Z(\mreg/_00093_ ) );
INV_X1 \mreg/_09671_ ( .A(\mreg/_04934_ ), .ZN(\mreg/_03705_ ) );
OR2_X1 \mreg/_09672_ ( .A1(\mreg/_03705_ ), .A2(\mreg/_04935_ ), .ZN(\mreg/_03706_ ) );
INV_X1 \mreg/_09673_ ( .A(\mreg/_03690_ ), .ZN(\mreg/_03707_ ) );
OR3_X1 \mreg/_09674_ ( .A1(\mreg/_03706_ ), .A2(\mreg/_03707_ ), .A3(\mreg/_04938_ ), .ZN(\mreg/_03708_ ) );
BUF_X4 \mreg/_09675_ ( .A(\mreg/_03695_ ), .Z(\mreg/_03709_ ) );
NOR2_X4 \mreg/_09676_ ( .A1(\mreg/_03708_ ), .A2(\mreg/_03709_ ), .ZN(\mreg/_03710_ ) );
BUF_X4 \mreg/_09677_ ( .A(\mreg/_03710_ ), .Z(\mreg/_03711_ ) );
MUX2_X1 \mreg/_09678_ ( .A(\mreg/_04262_ ), .B(\mreg/_04939_ ), .S(\mreg/_03711_ ), .Z(\mreg/_00094_ ) );
MUX2_X1 \mreg/_09679_ ( .A(\mreg/_04273_ ), .B(\mreg/_04950_ ), .S(\mreg/_03711_ ), .Z(\mreg/_00095_ ) );
MUX2_X1 \mreg/_09680_ ( .A(\mreg/_04284_ ), .B(\mreg/_04961_ ), .S(\mreg/_03711_ ), .Z(\mreg/_00096_ ) );
MUX2_X1 \mreg/_09681_ ( .A(\mreg/_04287_ ), .B(\mreg/_04964_ ), .S(\mreg/_03711_ ), .Z(\mreg/_00097_ ) );
MUX2_X1 \mreg/_09682_ ( .A(\mreg/_04288_ ), .B(\mreg/_04965_ ), .S(\mreg/_03711_ ), .Z(\mreg/_00098_ ) );
MUX2_X1 \mreg/_09683_ ( .A(\mreg/_04289_ ), .B(\mreg/_04966_ ), .S(\mreg/_03711_ ), .Z(\mreg/_00099_ ) );
MUX2_X1 \mreg/_09684_ ( .A(\mreg/_04290_ ), .B(\mreg/_04967_ ), .S(\mreg/_03711_ ), .Z(\mreg/_00100_ ) );
MUX2_X1 \mreg/_09685_ ( .A(\mreg/_04291_ ), .B(\mreg/_04968_ ), .S(\mreg/_03711_ ), .Z(\mreg/_00101_ ) );
MUX2_X1 \mreg/_09686_ ( .A(\mreg/_04292_ ), .B(\mreg/_04969_ ), .S(\mreg/_03711_ ), .Z(\mreg/_00102_ ) );
MUX2_X1 \mreg/_09687_ ( .A(\mreg/_04293_ ), .B(\mreg/_04970_ ), .S(\mreg/_03711_ ), .Z(\mreg/_00103_ ) );
BUF_X4 \mreg/_09688_ ( .A(\mreg/_03710_ ), .Z(\mreg/_03712_ ) );
MUX2_X1 \mreg/_09689_ ( .A(\mreg/_04263_ ), .B(\mreg/_04940_ ), .S(\mreg/_03712_ ), .Z(\mreg/_00104_ ) );
MUX2_X1 \mreg/_09690_ ( .A(\mreg/_04264_ ), .B(\mreg/_04941_ ), .S(\mreg/_03712_ ), .Z(\mreg/_00105_ ) );
MUX2_X1 \mreg/_09691_ ( .A(\mreg/_04265_ ), .B(\mreg/_04942_ ), .S(\mreg/_03712_ ), .Z(\mreg/_00106_ ) );
MUX2_X1 \mreg/_09692_ ( .A(\mreg/_04266_ ), .B(\mreg/_04943_ ), .S(\mreg/_03712_ ), .Z(\mreg/_00107_ ) );
MUX2_X1 \mreg/_09693_ ( .A(\mreg/_04267_ ), .B(\mreg/_04944_ ), .S(\mreg/_03712_ ), .Z(\mreg/_00108_ ) );
MUX2_X1 \mreg/_09694_ ( .A(\mreg/_04268_ ), .B(\mreg/_04945_ ), .S(\mreg/_03712_ ), .Z(\mreg/_00109_ ) );
MUX2_X1 \mreg/_09695_ ( .A(\mreg/_04269_ ), .B(\mreg/_04946_ ), .S(\mreg/_03712_ ), .Z(\mreg/_00110_ ) );
MUX2_X1 \mreg/_09696_ ( .A(\mreg/_04270_ ), .B(\mreg/_04947_ ), .S(\mreg/_03712_ ), .Z(\mreg/_00111_ ) );
MUX2_X1 \mreg/_09697_ ( .A(\mreg/_04271_ ), .B(\mreg/_04948_ ), .S(\mreg/_03712_ ), .Z(\mreg/_00112_ ) );
MUX2_X1 \mreg/_09698_ ( .A(\mreg/_04272_ ), .B(\mreg/_04949_ ), .S(\mreg/_03712_ ), .Z(\mreg/_00113_ ) );
BUF_X4 \mreg/_09699_ ( .A(\mreg/_03710_ ), .Z(\mreg/_03713_ ) );
MUX2_X1 \mreg/_09700_ ( .A(\mreg/_04274_ ), .B(\mreg/_04951_ ), .S(\mreg/_03713_ ), .Z(\mreg/_00114_ ) );
MUX2_X1 \mreg/_09701_ ( .A(\mreg/_04275_ ), .B(\mreg/_04952_ ), .S(\mreg/_03713_ ), .Z(\mreg/_00115_ ) );
MUX2_X1 \mreg/_09702_ ( .A(\mreg/_04276_ ), .B(\mreg/_04953_ ), .S(\mreg/_03713_ ), .Z(\mreg/_00116_ ) );
MUX2_X1 \mreg/_09703_ ( .A(\mreg/_04277_ ), .B(\mreg/_04954_ ), .S(\mreg/_03713_ ), .Z(\mreg/_00117_ ) );
MUX2_X1 \mreg/_09704_ ( .A(\mreg/_04278_ ), .B(\mreg/_04955_ ), .S(\mreg/_03713_ ), .Z(\mreg/_00118_ ) );
MUX2_X1 \mreg/_09705_ ( .A(\mreg/_04279_ ), .B(\mreg/_04956_ ), .S(\mreg/_03713_ ), .Z(\mreg/_00119_ ) );
MUX2_X1 \mreg/_09706_ ( .A(\mreg/_04280_ ), .B(\mreg/_04957_ ), .S(\mreg/_03713_ ), .Z(\mreg/_00120_ ) );
MUX2_X1 \mreg/_09707_ ( .A(\mreg/_04281_ ), .B(\mreg/_04958_ ), .S(\mreg/_03713_ ), .Z(\mreg/_00121_ ) );
MUX2_X1 \mreg/_09708_ ( .A(\mreg/_04282_ ), .B(\mreg/_04959_ ), .S(\mreg/_03713_ ), .Z(\mreg/_00122_ ) );
MUX2_X1 \mreg/_09709_ ( .A(\mreg/_04283_ ), .B(\mreg/_04960_ ), .S(\mreg/_03713_ ), .Z(\mreg/_00123_ ) );
MUX2_X1 \mreg/_09710_ ( .A(\mreg/_04285_ ), .B(\mreg/_04962_ ), .S(\mreg/_03710_ ), .Z(\mreg/_00124_ ) );
MUX2_X1 \mreg/_09711_ ( .A(\mreg/_04286_ ), .B(\mreg/_04963_ ), .S(\mreg/_03710_ ), .Z(\mreg/_00125_ ) );
BUF_X2 \mreg/_09712_ ( .A(\mreg/_03692_ ), .Z(\mreg/_03714_ ) );
NAND4_X1 \mreg/_09713_ ( .A1(\mreg/_03690_ ), .A2(\mreg/_03714_ ), .A3(\mreg/_03705_ ), .A4(\mreg/_04935_ ), .ZN(\mreg/_03715_ ) );
NOR2_X1 \mreg/_09714_ ( .A1(\mreg/_03696_ ), .A2(\mreg/_03715_ ), .ZN(\mreg/_03716_ ) );
BUF_X4 \mreg/_09715_ ( .A(\mreg/_03716_ ), .Z(\mreg/_03717_ ) );
MUX2_X1 \mreg/_09716_ ( .A(\mreg/_04614_ ), .B(\mreg/_04939_ ), .S(\mreg/_03717_ ), .Z(\mreg/_00126_ ) );
MUX2_X1 \mreg/_09717_ ( .A(\mreg/_04625_ ), .B(\mreg/_04950_ ), .S(\mreg/_03717_ ), .Z(\mreg/_00127_ ) );
MUX2_X1 \mreg/_09718_ ( .A(\mreg/_04636_ ), .B(\mreg/_04961_ ), .S(\mreg/_03717_ ), .Z(\mreg/_00128_ ) );
MUX2_X1 \mreg/_09719_ ( .A(\mreg/_04639_ ), .B(\mreg/_04964_ ), .S(\mreg/_03717_ ), .Z(\mreg/_00129_ ) );
MUX2_X1 \mreg/_09720_ ( .A(\mreg/_04640_ ), .B(\mreg/_04965_ ), .S(\mreg/_03717_ ), .Z(\mreg/_00130_ ) );
MUX2_X1 \mreg/_09721_ ( .A(\mreg/_04641_ ), .B(\mreg/_04966_ ), .S(\mreg/_03717_ ), .Z(\mreg/_00131_ ) );
MUX2_X1 \mreg/_09722_ ( .A(\mreg/_04642_ ), .B(\mreg/_04967_ ), .S(\mreg/_03717_ ), .Z(\mreg/_00132_ ) );
MUX2_X1 \mreg/_09723_ ( .A(\mreg/_04643_ ), .B(\mreg/_04968_ ), .S(\mreg/_03717_ ), .Z(\mreg/_00133_ ) );
MUX2_X1 \mreg/_09724_ ( .A(\mreg/_04644_ ), .B(\mreg/_04969_ ), .S(\mreg/_03717_ ), .Z(\mreg/_00134_ ) );
MUX2_X1 \mreg/_09725_ ( .A(\mreg/_04645_ ), .B(\mreg/_04970_ ), .S(\mreg/_03717_ ), .Z(\mreg/_00135_ ) );
BUF_X4 \mreg/_09726_ ( .A(\mreg/_03716_ ), .Z(\mreg/_03718_ ) );
MUX2_X1 \mreg/_09727_ ( .A(\mreg/_04615_ ), .B(\mreg/_04940_ ), .S(\mreg/_03718_ ), .Z(\mreg/_00136_ ) );
MUX2_X1 \mreg/_09728_ ( .A(\mreg/_04616_ ), .B(\mreg/_04941_ ), .S(\mreg/_03718_ ), .Z(\mreg/_00137_ ) );
MUX2_X1 \mreg/_09729_ ( .A(\mreg/_04617_ ), .B(\mreg/_04942_ ), .S(\mreg/_03718_ ), .Z(\mreg/_00138_ ) );
MUX2_X1 \mreg/_09730_ ( .A(\mreg/_04618_ ), .B(\mreg/_04943_ ), .S(\mreg/_03718_ ), .Z(\mreg/_00139_ ) );
MUX2_X1 \mreg/_09731_ ( .A(\mreg/_04619_ ), .B(\mreg/_04944_ ), .S(\mreg/_03718_ ), .Z(\mreg/_00140_ ) );
MUX2_X1 \mreg/_09732_ ( .A(\mreg/_04620_ ), .B(\mreg/_04945_ ), .S(\mreg/_03718_ ), .Z(\mreg/_00141_ ) );
MUX2_X1 \mreg/_09733_ ( .A(\mreg/_04621_ ), .B(\mreg/_04946_ ), .S(\mreg/_03718_ ), .Z(\mreg/_00142_ ) );
MUX2_X1 \mreg/_09734_ ( .A(\mreg/_04622_ ), .B(\mreg/_04947_ ), .S(\mreg/_03718_ ), .Z(\mreg/_00143_ ) );
MUX2_X1 \mreg/_09735_ ( .A(\mreg/_04623_ ), .B(\mreg/_04948_ ), .S(\mreg/_03718_ ), .Z(\mreg/_00144_ ) );
MUX2_X1 \mreg/_09736_ ( .A(\mreg/_04624_ ), .B(\mreg/_04949_ ), .S(\mreg/_03718_ ), .Z(\mreg/_00145_ ) );
BUF_X4 \mreg/_09737_ ( .A(\mreg/_03716_ ), .Z(\mreg/_03719_ ) );
MUX2_X1 \mreg/_09738_ ( .A(\mreg/_04626_ ), .B(\mreg/_04951_ ), .S(\mreg/_03719_ ), .Z(\mreg/_00146_ ) );
MUX2_X1 \mreg/_09739_ ( .A(\mreg/_04627_ ), .B(\mreg/_04952_ ), .S(\mreg/_03719_ ), .Z(\mreg/_00147_ ) );
MUX2_X1 \mreg/_09740_ ( .A(\mreg/_04628_ ), .B(\mreg/_04953_ ), .S(\mreg/_03719_ ), .Z(\mreg/_00148_ ) );
MUX2_X1 \mreg/_09741_ ( .A(\mreg/_04629_ ), .B(\mreg/_04954_ ), .S(\mreg/_03719_ ), .Z(\mreg/_00149_ ) );
MUX2_X1 \mreg/_09742_ ( .A(\mreg/_04630_ ), .B(\mreg/_04955_ ), .S(\mreg/_03719_ ), .Z(\mreg/_00150_ ) );
MUX2_X1 \mreg/_09743_ ( .A(\mreg/_04631_ ), .B(\mreg/_04956_ ), .S(\mreg/_03719_ ), .Z(\mreg/_00151_ ) );
MUX2_X1 \mreg/_09744_ ( .A(\mreg/_04632_ ), .B(\mreg/_04957_ ), .S(\mreg/_03719_ ), .Z(\mreg/_00152_ ) );
MUX2_X1 \mreg/_09745_ ( .A(\mreg/_04633_ ), .B(\mreg/_04958_ ), .S(\mreg/_03719_ ), .Z(\mreg/_00153_ ) );
MUX2_X1 \mreg/_09746_ ( .A(\mreg/_04634_ ), .B(\mreg/_04959_ ), .S(\mreg/_03719_ ), .Z(\mreg/_00154_ ) );
MUX2_X1 \mreg/_09747_ ( .A(\mreg/_04635_ ), .B(\mreg/_04960_ ), .S(\mreg/_03719_ ), .Z(\mreg/_00155_ ) );
MUX2_X1 \mreg/_09748_ ( .A(\mreg/_04637_ ), .B(\mreg/_04962_ ), .S(\mreg/_03716_ ), .Z(\mreg/_00156_ ) );
MUX2_X1 \mreg/_09749_ ( .A(\mreg/_04638_ ), .B(\mreg/_04963_ ), .S(\mreg/_03716_ ), .Z(\mreg/_00157_ ) );
NAND4_X1 \mreg/_09750_ ( .A1(\mreg/_03690_ ), .A2(\mreg/_03714_ ), .A3(\mreg/_04934_ ), .A4(\mreg/_04935_ ), .ZN(\mreg/_03720_ ) );
NOR2_X1 \mreg/_09751_ ( .A1(\mreg/_03696_ ), .A2(\mreg/_03720_ ), .ZN(\mreg/_03721_ ) );
BUF_X4 \mreg/_09752_ ( .A(\mreg/_03721_ ), .Z(\mreg/_03722_ ) );
MUX2_X1 \mreg/_09753_ ( .A(\mreg/_04710_ ), .B(\mreg/_04939_ ), .S(\mreg/_03722_ ), .Z(\mreg/_00158_ ) );
MUX2_X1 \mreg/_09754_ ( .A(\mreg/_04721_ ), .B(\mreg/_04950_ ), .S(\mreg/_03722_ ), .Z(\mreg/_00159_ ) );
MUX2_X1 \mreg/_09755_ ( .A(\mreg/_04732_ ), .B(\mreg/_04961_ ), .S(\mreg/_03722_ ), .Z(\mreg/_00160_ ) );
MUX2_X1 \mreg/_09756_ ( .A(\mreg/_04735_ ), .B(\mreg/_04964_ ), .S(\mreg/_03722_ ), .Z(\mreg/_00161_ ) );
MUX2_X1 \mreg/_09757_ ( .A(\mreg/_04736_ ), .B(\mreg/_04965_ ), .S(\mreg/_03722_ ), .Z(\mreg/_00162_ ) );
MUX2_X1 \mreg/_09758_ ( .A(\mreg/_04737_ ), .B(\mreg/_04966_ ), .S(\mreg/_03722_ ), .Z(\mreg/_00163_ ) );
MUX2_X1 \mreg/_09759_ ( .A(\mreg/_04738_ ), .B(\mreg/_04967_ ), .S(\mreg/_03722_ ), .Z(\mreg/_00164_ ) );
MUX2_X1 \mreg/_09760_ ( .A(\mreg/_04739_ ), .B(\mreg/_04968_ ), .S(\mreg/_03722_ ), .Z(\mreg/_00165_ ) );
MUX2_X1 \mreg/_09761_ ( .A(\mreg/_04740_ ), .B(\mreg/_04969_ ), .S(\mreg/_03722_ ), .Z(\mreg/_00166_ ) );
MUX2_X1 \mreg/_09762_ ( .A(\mreg/_04741_ ), .B(\mreg/_04970_ ), .S(\mreg/_03722_ ), .Z(\mreg/_00167_ ) );
BUF_X4 \mreg/_09763_ ( .A(\mreg/_03721_ ), .Z(\mreg/_03723_ ) );
MUX2_X1 \mreg/_09764_ ( .A(\mreg/_04711_ ), .B(\mreg/_04940_ ), .S(\mreg/_03723_ ), .Z(\mreg/_00168_ ) );
MUX2_X1 \mreg/_09765_ ( .A(\mreg/_04712_ ), .B(\mreg/_04941_ ), .S(\mreg/_03723_ ), .Z(\mreg/_00169_ ) );
MUX2_X1 \mreg/_09766_ ( .A(\mreg/_04713_ ), .B(\mreg/_04942_ ), .S(\mreg/_03723_ ), .Z(\mreg/_00170_ ) );
MUX2_X1 \mreg/_09767_ ( .A(\mreg/_04714_ ), .B(\mreg/_04943_ ), .S(\mreg/_03723_ ), .Z(\mreg/_00171_ ) );
MUX2_X1 \mreg/_09768_ ( .A(\mreg/_04715_ ), .B(\mreg/_04944_ ), .S(\mreg/_03723_ ), .Z(\mreg/_00172_ ) );
MUX2_X1 \mreg/_09769_ ( .A(\mreg/_04716_ ), .B(\mreg/_04945_ ), .S(\mreg/_03723_ ), .Z(\mreg/_00173_ ) );
MUX2_X1 \mreg/_09770_ ( .A(\mreg/_04717_ ), .B(\mreg/_04946_ ), .S(\mreg/_03723_ ), .Z(\mreg/_00174_ ) );
MUX2_X1 \mreg/_09771_ ( .A(\mreg/_04718_ ), .B(\mreg/_04947_ ), .S(\mreg/_03723_ ), .Z(\mreg/_00175_ ) );
MUX2_X1 \mreg/_09772_ ( .A(\mreg/_04719_ ), .B(\mreg/_04948_ ), .S(\mreg/_03723_ ), .Z(\mreg/_00176_ ) );
MUX2_X1 \mreg/_09773_ ( .A(\mreg/_04720_ ), .B(\mreg/_04949_ ), .S(\mreg/_03723_ ), .Z(\mreg/_00177_ ) );
BUF_X4 \mreg/_09774_ ( .A(\mreg/_03721_ ), .Z(\mreg/_03724_ ) );
MUX2_X1 \mreg/_09775_ ( .A(\mreg/_04722_ ), .B(\mreg/_04951_ ), .S(\mreg/_03724_ ), .Z(\mreg/_00178_ ) );
MUX2_X1 \mreg/_09776_ ( .A(\mreg/_04723_ ), .B(\mreg/_04952_ ), .S(\mreg/_03724_ ), .Z(\mreg/_00179_ ) );
MUX2_X1 \mreg/_09777_ ( .A(\mreg/_04724_ ), .B(\mreg/_04953_ ), .S(\mreg/_03724_ ), .Z(\mreg/_00180_ ) );
MUX2_X1 \mreg/_09778_ ( .A(\mreg/_04725_ ), .B(\mreg/_04954_ ), .S(\mreg/_03724_ ), .Z(\mreg/_00181_ ) );
MUX2_X1 \mreg/_09779_ ( .A(\mreg/_04726_ ), .B(\mreg/_04955_ ), .S(\mreg/_03724_ ), .Z(\mreg/_00182_ ) );
MUX2_X1 \mreg/_09780_ ( .A(\mreg/_04727_ ), .B(\mreg/_04956_ ), .S(\mreg/_03724_ ), .Z(\mreg/_00183_ ) );
MUX2_X1 \mreg/_09781_ ( .A(\mreg/_04728_ ), .B(\mreg/_04957_ ), .S(\mreg/_03724_ ), .Z(\mreg/_00184_ ) );
MUX2_X1 \mreg/_09782_ ( .A(\mreg/_04729_ ), .B(\mreg/_04958_ ), .S(\mreg/_03724_ ), .Z(\mreg/_00185_ ) );
MUX2_X1 \mreg/_09783_ ( .A(\mreg/_04730_ ), .B(\mreg/_04959_ ), .S(\mreg/_03724_ ), .Z(\mreg/_00186_ ) );
MUX2_X1 \mreg/_09784_ ( .A(\mreg/_04731_ ), .B(\mreg/_04960_ ), .S(\mreg/_03724_ ), .Z(\mreg/_00187_ ) );
MUX2_X1 \mreg/_09785_ ( .A(\mreg/_04733_ ), .B(\mreg/_04962_ ), .S(\mreg/_03721_ ), .Z(\mreg/_00188_ ) );
MUX2_X1 \mreg/_09786_ ( .A(\mreg/_04734_ ), .B(\mreg/_04963_ ), .S(\mreg/_03721_ ), .Z(\mreg/_00189_ ) );
INV_X1 \mreg/_09787_ ( .A(\mreg/_04936_ ), .ZN(\mreg/_03725_ ) );
OR2_X1 \mreg/_09788_ ( .A1(\mreg/_03725_ ), .A2(\mreg/_04937_ ), .ZN(\mreg/_03726_ ) );
INV_X1 \mreg/_09789_ ( .A(\mreg/_03691_ ), .ZN(\mreg/_03727_ ) );
OR3_X1 \mreg/_09790_ ( .A1(\mreg/_03726_ ), .A2(\mreg/_03727_ ), .A3(\mreg/_04938_ ), .ZN(\mreg/_03728_ ) );
NOR2_X4 \mreg/_09791_ ( .A1(\mreg/_03728_ ), .A2(\mreg/_03709_ ), .ZN(\mreg/_03729_ ) );
BUF_X4 \mreg/_09792_ ( .A(\mreg/_03729_ ), .Z(\mreg/_03730_ ) );
MUX2_X1 \mreg/_09793_ ( .A(\mreg/_04742_ ), .B(\mreg/_04939_ ), .S(\mreg/_03730_ ), .Z(\mreg/_00190_ ) );
MUX2_X1 \mreg/_09794_ ( .A(\mreg/_04753_ ), .B(\mreg/_04950_ ), .S(\mreg/_03730_ ), .Z(\mreg/_00191_ ) );
MUX2_X1 \mreg/_09795_ ( .A(\mreg/_04764_ ), .B(\mreg/_04961_ ), .S(\mreg/_03730_ ), .Z(\mreg/_00192_ ) );
MUX2_X1 \mreg/_09796_ ( .A(\mreg/_04767_ ), .B(\mreg/_04964_ ), .S(\mreg/_03730_ ), .Z(\mreg/_00193_ ) );
MUX2_X1 \mreg/_09797_ ( .A(\mreg/_04768_ ), .B(\mreg/_04965_ ), .S(\mreg/_03730_ ), .Z(\mreg/_00194_ ) );
MUX2_X1 \mreg/_09798_ ( .A(\mreg/_04769_ ), .B(\mreg/_04966_ ), .S(\mreg/_03730_ ), .Z(\mreg/_00195_ ) );
MUX2_X1 \mreg/_09799_ ( .A(\mreg/_04770_ ), .B(\mreg/_04967_ ), .S(\mreg/_03730_ ), .Z(\mreg/_00196_ ) );
MUX2_X1 \mreg/_09800_ ( .A(\mreg/_04771_ ), .B(\mreg/_04968_ ), .S(\mreg/_03730_ ), .Z(\mreg/_00197_ ) );
MUX2_X1 \mreg/_09801_ ( .A(\mreg/_04772_ ), .B(\mreg/_04969_ ), .S(\mreg/_03730_ ), .Z(\mreg/_00198_ ) );
MUX2_X1 \mreg/_09802_ ( .A(\mreg/_04773_ ), .B(\mreg/_04970_ ), .S(\mreg/_03730_ ), .Z(\mreg/_00199_ ) );
BUF_X4 \mreg/_09803_ ( .A(\mreg/_03729_ ), .Z(\mreg/_03731_ ) );
MUX2_X1 \mreg/_09804_ ( .A(\mreg/_04743_ ), .B(\mreg/_04940_ ), .S(\mreg/_03731_ ), .Z(\mreg/_00200_ ) );
MUX2_X1 \mreg/_09805_ ( .A(\mreg/_04744_ ), .B(\mreg/_04941_ ), .S(\mreg/_03731_ ), .Z(\mreg/_00201_ ) );
MUX2_X1 \mreg/_09806_ ( .A(\mreg/_04745_ ), .B(\mreg/_04942_ ), .S(\mreg/_03731_ ), .Z(\mreg/_00202_ ) );
MUX2_X1 \mreg/_09807_ ( .A(\mreg/_04746_ ), .B(\mreg/_04943_ ), .S(\mreg/_03731_ ), .Z(\mreg/_00203_ ) );
MUX2_X1 \mreg/_09808_ ( .A(\mreg/_04747_ ), .B(\mreg/_04944_ ), .S(\mreg/_03731_ ), .Z(\mreg/_00204_ ) );
MUX2_X1 \mreg/_09809_ ( .A(\mreg/_04748_ ), .B(\mreg/_04945_ ), .S(\mreg/_03731_ ), .Z(\mreg/_00205_ ) );
MUX2_X1 \mreg/_09810_ ( .A(\mreg/_04749_ ), .B(\mreg/_04946_ ), .S(\mreg/_03731_ ), .Z(\mreg/_00206_ ) );
MUX2_X1 \mreg/_09811_ ( .A(\mreg/_04750_ ), .B(\mreg/_04947_ ), .S(\mreg/_03731_ ), .Z(\mreg/_00207_ ) );
MUX2_X1 \mreg/_09812_ ( .A(\mreg/_04751_ ), .B(\mreg/_04948_ ), .S(\mreg/_03731_ ), .Z(\mreg/_00208_ ) );
MUX2_X1 \mreg/_09813_ ( .A(\mreg/_04752_ ), .B(\mreg/_04949_ ), .S(\mreg/_03731_ ), .Z(\mreg/_00209_ ) );
BUF_X4 \mreg/_09814_ ( .A(\mreg/_03729_ ), .Z(\mreg/_03732_ ) );
MUX2_X1 \mreg/_09815_ ( .A(\mreg/_04754_ ), .B(\mreg/_04951_ ), .S(\mreg/_03732_ ), .Z(\mreg/_00210_ ) );
MUX2_X1 \mreg/_09816_ ( .A(\mreg/_04755_ ), .B(\mreg/_04952_ ), .S(\mreg/_03732_ ), .Z(\mreg/_00211_ ) );
MUX2_X1 \mreg/_09817_ ( .A(\mreg/_04756_ ), .B(\mreg/_04953_ ), .S(\mreg/_03732_ ), .Z(\mreg/_00212_ ) );
MUX2_X1 \mreg/_09818_ ( .A(\mreg/_04757_ ), .B(\mreg/_04954_ ), .S(\mreg/_03732_ ), .Z(\mreg/_00213_ ) );
MUX2_X1 \mreg/_09819_ ( .A(\mreg/_04758_ ), .B(\mreg/_04955_ ), .S(\mreg/_03732_ ), .Z(\mreg/_00214_ ) );
MUX2_X1 \mreg/_09820_ ( .A(\mreg/_04759_ ), .B(\mreg/_04956_ ), .S(\mreg/_03732_ ), .Z(\mreg/_00215_ ) );
MUX2_X1 \mreg/_09821_ ( .A(\mreg/_04760_ ), .B(\mreg/_04957_ ), .S(\mreg/_03732_ ), .Z(\mreg/_00216_ ) );
MUX2_X1 \mreg/_09822_ ( .A(\mreg/_04761_ ), .B(\mreg/_04958_ ), .S(\mreg/_03732_ ), .Z(\mreg/_00217_ ) );
MUX2_X1 \mreg/_09823_ ( .A(\mreg/_04762_ ), .B(\mreg/_04959_ ), .S(\mreg/_03732_ ), .Z(\mreg/_00218_ ) );
MUX2_X1 \mreg/_09824_ ( .A(\mreg/_04763_ ), .B(\mreg/_04960_ ), .S(\mreg/_03732_ ), .Z(\mreg/_00219_ ) );
MUX2_X1 \mreg/_09825_ ( .A(\mreg/_04765_ ), .B(\mreg/_04962_ ), .S(\mreg/_03729_ ), .Z(\mreg/_00220_ ) );
MUX2_X1 \mreg/_09826_ ( .A(\mreg/_04766_ ), .B(\mreg/_04963_ ), .S(\mreg/_03729_ ), .Z(\mreg/_00221_ ) );
NOR2_X1 \mreg/_09827_ ( .A1(\mreg/_03706_ ), .A2(\mreg/_03726_ ), .ZN(\mreg/_03733_ ) );
NAND2_X1 \mreg/_09828_ ( .A1(\mreg/_03733_ ), .A2(\mreg/_03714_ ), .ZN(\mreg/_03734_ ) );
NOR2_X1 \mreg/_09829_ ( .A1(\mreg/_03734_ ), .A2(\mreg/_03709_ ), .ZN(\mreg/_03735_ ) );
BUF_X4 \mreg/_09830_ ( .A(\mreg/_03735_ ), .Z(\mreg/_03736_ ) );
MUX2_X1 \mreg/_09831_ ( .A(\mreg/_04774_ ), .B(\mreg/_04939_ ), .S(\mreg/_03736_ ), .Z(\mreg/_00222_ ) );
MUX2_X1 \mreg/_09832_ ( .A(\mreg/_04785_ ), .B(\mreg/_04950_ ), .S(\mreg/_03736_ ), .Z(\mreg/_00223_ ) );
MUX2_X1 \mreg/_09833_ ( .A(\mreg/_04796_ ), .B(\mreg/_04961_ ), .S(\mreg/_03736_ ), .Z(\mreg/_00224_ ) );
MUX2_X1 \mreg/_09834_ ( .A(\mreg/_04799_ ), .B(\mreg/_04964_ ), .S(\mreg/_03736_ ), .Z(\mreg/_00225_ ) );
MUX2_X1 \mreg/_09835_ ( .A(\mreg/_04800_ ), .B(\mreg/_04965_ ), .S(\mreg/_03736_ ), .Z(\mreg/_00226_ ) );
MUX2_X1 \mreg/_09836_ ( .A(\mreg/_04801_ ), .B(\mreg/_04966_ ), .S(\mreg/_03736_ ), .Z(\mreg/_00227_ ) );
MUX2_X1 \mreg/_09837_ ( .A(\mreg/_04802_ ), .B(\mreg/_04967_ ), .S(\mreg/_03736_ ), .Z(\mreg/_00228_ ) );
MUX2_X1 \mreg/_09838_ ( .A(\mreg/_04803_ ), .B(\mreg/_04968_ ), .S(\mreg/_03736_ ), .Z(\mreg/_00229_ ) );
MUX2_X1 \mreg/_09839_ ( .A(\mreg/_04804_ ), .B(\mreg/_04969_ ), .S(\mreg/_03736_ ), .Z(\mreg/_00230_ ) );
MUX2_X1 \mreg/_09840_ ( .A(\mreg/_04805_ ), .B(\mreg/_04970_ ), .S(\mreg/_03736_ ), .Z(\mreg/_00231_ ) );
BUF_X4 \mreg/_09841_ ( .A(\mreg/_03735_ ), .Z(\mreg/_03737_ ) );
MUX2_X1 \mreg/_09842_ ( .A(\mreg/_04775_ ), .B(\mreg/_04940_ ), .S(\mreg/_03737_ ), .Z(\mreg/_00232_ ) );
MUX2_X1 \mreg/_09843_ ( .A(\mreg/_04776_ ), .B(\mreg/_04941_ ), .S(\mreg/_03737_ ), .Z(\mreg/_00233_ ) );
MUX2_X1 \mreg/_09844_ ( .A(\mreg/_04777_ ), .B(\mreg/_04942_ ), .S(\mreg/_03737_ ), .Z(\mreg/_00234_ ) );
MUX2_X1 \mreg/_09845_ ( .A(\mreg/_04778_ ), .B(\mreg/_04943_ ), .S(\mreg/_03737_ ), .Z(\mreg/_00235_ ) );
MUX2_X1 \mreg/_09846_ ( .A(\mreg/_04779_ ), .B(\mreg/_04944_ ), .S(\mreg/_03737_ ), .Z(\mreg/_00236_ ) );
MUX2_X1 \mreg/_09847_ ( .A(\mreg/_04780_ ), .B(\mreg/_04945_ ), .S(\mreg/_03737_ ), .Z(\mreg/_00237_ ) );
MUX2_X1 \mreg/_09848_ ( .A(\mreg/_04781_ ), .B(\mreg/_04946_ ), .S(\mreg/_03737_ ), .Z(\mreg/_00238_ ) );
MUX2_X1 \mreg/_09849_ ( .A(\mreg/_04782_ ), .B(\mreg/_04947_ ), .S(\mreg/_03737_ ), .Z(\mreg/_00239_ ) );
MUX2_X1 \mreg/_09850_ ( .A(\mreg/_04783_ ), .B(\mreg/_04948_ ), .S(\mreg/_03737_ ), .Z(\mreg/_00240_ ) );
MUX2_X1 \mreg/_09851_ ( .A(\mreg/_04784_ ), .B(\mreg/_04949_ ), .S(\mreg/_03737_ ), .Z(\mreg/_00241_ ) );
BUF_X4 \mreg/_09852_ ( .A(\mreg/_03735_ ), .Z(\mreg/_03738_ ) );
MUX2_X1 \mreg/_09853_ ( .A(\mreg/_04786_ ), .B(\mreg/_04951_ ), .S(\mreg/_03738_ ), .Z(\mreg/_00242_ ) );
MUX2_X1 \mreg/_09854_ ( .A(\mreg/_04787_ ), .B(\mreg/_04952_ ), .S(\mreg/_03738_ ), .Z(\mreg/_00243_ ) );
MUX2_X1 \mreg/_09855_ ( .A(\mreg/_04788_ ), .B(\mreg/_04953_ ), .S(\mreg/_03738_ ), .Z(\mreg/_00244_ ) );
MUX2_X1 \mreg/_09856_ ( .A(\mreg/_04789_ ), .B(\mreg/_04954_ ), .S(\mreg/_03738_ ), .Z(\mreg/_00245_ ) );
MUX2_X1 \mreg/_09857_ ( .A(\mreg/_04790_ ), .B(\mreg/_04955_ ), .S(\mreg/_03738_ ), .Z(\mreg/_00246_ ) );
MUX2_X1 \mreg/_09858_ ( .A(\mreg/_04791_ ), .B(\mreg/_04956_ ), .S(\mreg/_03738_ ), .Z(\mreg/_00247_ ) );
MUX2_X1 \mreg/_09859_ ( .A(\mreg/_04792_ ), .B(\mreg/_04957_ ), .S(\mreg/_03738_ ), .Z(\mreg/_00248_ ) );
MUX2_X1 \mreg/_09860_ ( .A(\mreg/_04793_ ), .B(\mreg/_04958_ ), .S(\mreg/_03738_ ), .Z(\mreg/_00249_ ) );
MUX2_X1 \mreg/_09861_ ( .A(\mreg/_04794_ ), .B(\mreg/_04959_ ), .S(\mreg/_03738_ ), .Z(\mreg/_00250_ ) );
MUX2_X1 \mreg/_09862_ ( .A(\mreg/_04795_ ), .B(\mreg/_04960_ ), .S(\mreg/_03738_ ), .Z(\mreg/_00251_ ) );
MUX2_X1 \mreg/_09863_ ( .A(\mreg/_04797_ ), .B(\mreg/_04962_ ), .S(\mreg/_03735_ ), .Z(\mreg/_00252_ ) );
MUX2_X1 \mreg/_09864_ ( .A(\mreg/_04798_ ), .B(\mreg/_04963_ ), .S(\mreg/_03735_ ), .Z(\mreg/_00253_ ) );
NAND2_X1 \mreg/_09865_ ( .A1(\mreg/_03705_ ), .A2(\mreg/_04935_ ), .ZN(\mreg/_03739_ ) );
OR3_X1 \mreg/_09866_ ( .A1(\mreg/_03726_ ), .A2(\mreg/_04938_ ), .A3(\mreg/_03739_ ), .ZN(\mreg/_03740_ ) );
NOR2_X1 \mreg/_09867_ ( .A1(\mreg/_03740_ ), .A2(\mreg/_03709_ ), .ZN(\mreg/_03741_ ) );
BUF_X4 \mreg/_09868_ ( .A(\mreg/_03741_ ), .Z(\mreg/_03742_ ) );
MUX2_X1 \mreg/_09869_ ( .A(\mreg/_04806_ ), .B(\mreg/_04939_ ), .S(\mreg/_03742_ ), .Z(\mreg/_00254_ ) );
MUX2_X1 \mreg/_09870_ ( .A(\mreg/_04817_ ), .B(\mreg/_04950_ ), .S(\mreg/_03742_ ), .Z(\mreg/_00255_ ) );
MUX2_X1 \mreg/_09871_ ( .A(\mreg/_04828_ ), .B(\mreg/_04961_ ), .S(\mreg/_03742_ ), .Z(\mreg/_00256_ ) );
MUX2_X1 \mreg/_09872_ ( .A(\mreg/_04831_ ), .B(\mreg/_04964_ ), .S(\mreg/_03742_ ), .Z(\mreg/_00257_ ) );
MUX2_X1 \mreg/_09873_ ( .A(\mreg/_04832_ ), .B(\mreg/_04965_ ), .S(\mreg/_03742_ ), .Z(\mreg/_00258_ ) );
MUX2_X1 \mreg/_09874_ ( .A(\mreg/_04833_ ), .B(\mreg/_04966_ ), .S(\mreg/_03742_ ), .Z(\mreg/_00259_ ) );
MUX2_X1 \mreg/_09875_ ( .A(\mreg/_04834_ ), .B(\mreg/_04967_ ), .S(\mreg/_03742_ ), .Z(\mreg/_00260_ ) );
MUX2_X1 \mreg/_09876_ ( .A(\mreg/_04835_ ), .B(\mreg/_04968_ ), .S(\mreg/_03742_ ), .Z(\mreg/_00261_ ) );
MUX2_X1 \mreg/_09877_ ( .A(\mreg/_04836_ ), .B(\mreg/_04969_ ), .S(\mreg/_03742_ ), .Z(\mreg/_00262_ ) );
MUX2_X1 \mreg/_09878_ ( .A(\mreg/_04837_ ), .B(\mreg/_04970_ ), .S(\mreg/_03742_ ), .Z(\mreg/_00263_ ) );
BUF_X4 \mreg/_09879_ ( .A(\mreg/_03741_ ), .Z(\mreg/_03743_ ) );
MUX2_X1 \mreg/_09880_ ( .A(\mreg/_04807_ ), .B(\mreg/_04940_ ), .S(\mreg/_03743_ ), .Z(\mreg/_00264_ ) );
MUX2_X1 \mreg/_09881_ ( .A(\mreg/_04808_ ), .B(\mreg/_04941_ ), .S(\mreg/_03743_ ), .Z(\mreg/_00265_ ) );
MUX2_X1 \mreg/_09882_ ( .A(\mreg/_04809_ ), .B(\mreg/_04942_ ), .S(\mreg/_03743_ ), .Z(\mreg/_00266_ ) );
MUX2_X1 \mreg/_09883_ ( .A(\mreg/_04810_ ), .B(\mreg/_04943_ ), .S(\mreg/_03743_ ), .Z(\mreg/_00267_ ) );
MUX2_X1 \mreg/_09884_ ( .A(\mreg/_04811_ ), .B(\mreg/_04944_ ), .S(\mreg/_03743_ ), .Z(\mreg/_00268_ ) );
MUX2_X1 \mreg/_09885_ ( .A(\mreg/_04812_ ), .B(\mreg/_04945_ ), .S(\mreg/_03743_ ), .Z(\mreg/_00269_ ) );
MUX2_X1 \mreg/_09886_ ( .A(\mreg/_04813_ ), .B(\mreg/_04946_ ), .S(\mreg/_03743_ ), .Z(\mreg/_00270_ ) );
MUX2_X1 \mreg/_09887_ ( .A(\mreg/_04814_ ), .B(\mreg/_04947_ ), .S(\mreg/_03743_ ), .Z(\mreg/_00271_ ) );
MUX2_X1 \mreg/_09888_ ( .A(\mreg/_04815_ ), .B(\mreg/_04948_ ), .S(\mreg/_03743_ ), .Z(\mreg/_00272_ ) );
MUX2_X1 \mreg/_09889_ ( .A(\mreg/_04816_ ), .B(\mreg/_04949_ ), .S(\mreg/_03743_ ), .Z(\mreg/_00273_ ) );
BUF_X4 \mreg/_09890_ ( .A(\mreg/_03741_ ), .Z(\mreg/_03744_ ) );
MUX2_X1 \mreg/_09891_ ( .A(\mreg/_04818_ ), .B(\mreg/_04951_ ), .S(\mreg/_03744_ ), .Z(\mreg/_00274_ ) );
MUX2_X1 \mreg/_09892_ ( .A(\mreg/_04819_ ), .B(\mreg/_04952_ ), .S(\mreg/_03744_ ), .Z(\mreg/_00275_ ) );
MUX2_X1 \mreg/_09893_ ( .A(\mreg/_04820_ ), .B(\mreg/_04953_ ), .S(\mreg/_03744_ ), .Z(\mreg/_00276_ ) );
MUX2_X1 \mreg/_09894_ ( .A(\mreg/_04821_ ), .B(\mreg/_04954_ ), .S(\mreg/_03744_ ), .Z(\mreg/_00277_ ) );
MUX2_X1 \mreg/_09895_ ( .A(\mreg/_04822_ ), .B(\mreg/_04955_ ), .S(\mreg/_03744_ ), .Z(\mreg/_00278_ ) );
MUX2_X1 \mreg/_09896_ ( .A(\mreg/_04823_ ), .B(\mreg/_04956_ ), .S(\mreg/_03744_ ), .Z(\mreg/_00279_ ) );
MUX2_X1 \mreg/_09897_ ( .A(\mreg/_04824_ ), .B(\mreg/_04957_ ), .S(\mreg/_03744_ ), .Z(\mreg/_00280_ ) );
MUX2_X1 \mreg/_09898_ ( .A(\mreg/_04825_ ), .B(\mreg/_04958_ ), .S(\mreg/_03744_ ), .Z(\mreg/_00281_ ) );
MUX2_X1 \mreg/_09899_ ( .A(\mreg/_04826_ ), .B(\mreg/_04959_ ), .S(\mreg/_03744_ ), .Z(\mreg/_00282_ ) );
MUX2_X1 \mreg/_09900_ ( .A(\mreg/_04827_ ), .B(\mreg/_04960_ ), .S(\mreg/_03744_ ), .Z(\mreg/_00283_ ) );
MUX2_X1 \mreg/_09901_ ( .A(\mreg/_04829_ ), .B(\mreg/_04962_ ), .S(\mreg/_03741_ ), .Z(\mreg/_00284_ ) );
MUX2_X1 \mreg/_09902_ ( .A(\mreg/_04830_ ), .B(\mreg/_04963_ ), .S(\mreg/_03741_ ), .Z(\mreg/_00285_ ) );
OR4_X1 \mreg/_09903_ ( .A1(\mreg/_04938_ ), .A2(\mreg/_03698_ ), .A3(\mreg/_03725_ ), .A4(\mreg/_04937_ ), .ZN(\mreg/_03745_ ) );
NOR2_X1 \mreg/_09904_ ( .A1(\mreg/_03745_ ), .A2(\mreg/_03709_ ), .ZN(\mreg/_03746_ ) );
BUF_X4 \mreg/_09905_ ( .A(\mreg/_03746_ ), .Z(\mreg/_03747_ ) );
MUX2_X1 \mreg/_09906_ ( .A(\mreg/_04838_ ), .B(\mreg/_04939_ ), .S(\mreg/_03747_ ), .Z(\mreg/_00286_ ) );
MUX2_X1 \mreg/_09907_ ( .A(\mreg/_04849_ ), .B(\mreg/_04950_ ), .S(\mreg/_03747_ ), .Z(\mreg/_00287_ ) );
MUX2_X1 \mreg/_09908_ ( .A(\mreg/_04860_ ), .B(\mreg/_04961_ ), .S(\mreg/_03747_ ), .Z(\mreg/_00288_ ) );
MUX2_X1 \mreg/_09909_ ( .A(\mreg/_04863_ ), .B(\mreg/_04964_ ), .S(\mreg/_03747_ ), .Z(\mreg/_00289_ ) );
MUX2_X1 \mreg/_09910_ ( .A(\mreg/_04864_ ), .B(\mreg/_04965_ ), .S(\mreg/_03747_ ), .Z(\mreg/_00290_ ) );
MUX2_X1 \mreg/_09911_ ( .A(\mreg/_04865_ ), .B(\mreg/_04966_ ), .S(\mreg/_03747_ ), .Z(\mreg/_00291_ ) );
MUX2_X1 \mreg/_09912_ ( .A(\mreg/_04866_ ), .B(\mreg/_04967_ ), .S(\mreg/_03747_ ), .Z(\mreg/_00292_ ) );
MUX2_X1 \mreg/_09913_ ( .A(\mreg/_04867_ ), .B(\mreg/_04968_ ), .S(\mreg/_03747_ ), .Z(\mreg/_00293_ ) );
MUX2_X1 \mreg/_09914_ ( .A(\mreg/_04868_ ), .B(\mreg/_04969_ ), .S(\mreg/_03747_ ), .Z(\mreg/_00294_ ) );
MUX2_X1 \mreg/_09915_ ( .A(\mreg/_04869_ ), .B(\mreg/_04970_ ), .S(\mreg/_03747_ ), .Z(\mreg/_00295_ ) );
BUF_X4 \mreg/_09916_ ( .A(\mreg/_03746_ ), .Z(\mreg/_03748_ ) );
MUX2_X1 \mreg/_09917_ ( .A(\mreg/_04839_ ), .B(\mreg/_04940_ ), .S(\mreg/_03748_ ), .Z(\mreg/_00296_ ) );
MUX2_X1 \mreg/_09918_ ( .A(\mreg/_04840_ ), .B(\mreg/_04941_ ), .S(\mreg/_03748_ ), .Z(\mreg/_00297_ ) );
MUX2_X1 \mreg/_09919_ ( .A(\mreg/_04841_ ), .B(\mreg/_04942_ ), .S(\mreg/_03748_ ), .Z(\mreg/_00298_ ) );
MUX2_X1 \mreg/_09920_ ( .A(\mreg/_04842_ ), .B(\mreg/_04943_ ), .S(\mreg/_03748_ ), .Z(\mreg/_00299_ ) );
MUX2_X1 \mreg/_09921_ ( .A(\mreg/_04843_ ), .B(\mreg/_04944_ ), .S(\mreg/_03748_ ), .Z(\mreg/_00300_ ) );
MUX2_X1 \mreg/_09922_ ( .A(\mreg/_04844_ ), .B(\mreg/_04945_ ), .S(\mreg/_03748_ ), .Z(\mreg/_00301_ ) );
MUX2_X1 \mreg/_09923_ ( .A(\mreg/_04845_ ), .B(\mreg/_04946_ ), .S(\mreg/_03748_ ), .Z(\mreg/_00302_ ) );
MUX2_X1 \mreg/_09924_ ( .A(\mreg/_04846_ ), .B(\mreg/_04947_ ), .S(\mreg/_03748_ ), .Z(\mreg/_00303_ ) );
MUX2_X1 \mreg/_09925_ ( .A(\mreg/_04847_ ), .B(\mreg/_04948_ ), .S(\mreg/_03748_ ), .Z(\mreg/_00304_ ) );
MUX2_X1 \mreg/_09926_ ( .A(\mreg/_04848_ ), .B(\mreg/_04949_ ), .S(\mreg/_03748_ ), .Z(\mreg/_00305_ ) );
BUF_X4 \mreg/_09927_ ( .A(\mreg/_03746_ ), .Z(\mreg/_03749_ ) );
MUX2_X1 \mreg/_09928_ ( .A(\mreg/_04850_ ), .B(\mreg/_04951_ ), .S(\mreg/_03749_ ), .Z(\mreg/_00306_ ) );
MUX2_X1 \mreg/_09929_ ( .A(\mreg/_04851_ ), .B(\mreg/_04952_ ), .S(\mreg/_03749_ ), .Z(\mreg/_00307_ ) );
MUX2_X1 \mreg/_09930_ ( .A(\mreg/_04852_ ), .B(\mreg/_04953_ ), .S(\mreg/_03749_ ), .Z(\mreg/_00308_ ) );
MUX2_X1 \mreg/_09931_ ( .A(\mreg/_04853_ ), .B(\mreg/_04954_ ), .S(\mreg/_03749_ ), .Z(\mreg/_00309_ ) );
MUX2_X1 \mreg/_09932_ ( .A(\mreg/_04854_ ), .B(\mreg/_04955_ ), .S(\mreg/_03749_ ), .Z(\mreg/_00310_ ) );
MUX2_X1 \mreg/_09933_ ( .A(\mreg/_04855_ ), .B(\mreg/_04956_ ), .S(\mreg/_03749_ ), .Z(\mreg/_00311_ ) );
MUX2_X1 \mreg/_09934_ ( .A(\mreg/_04856_ ), .B(\mreg/_04957_ ), .S(\mreg/_03749_ ), .Z(\mreg/_00312_ ) );
MUX2_X1 \mreg/_09935_ ( .A(\mreg/_04857_ ), .B(\mreg/_04958_ ), .S(\mreg/_03749_ ), .Z(\mreg/_00313_ ) );
MUX2_X1 \mreg/_09936_ ( .A(\mreg/_04858_ ), .B(\mreg/_04959_ ), .S(\mreg/_03749_ ), .Z(\mreg/_00314_ ) );
MUX2_X1 \mreg/_09937_ ( .A(\mreg/_04859_ ), .B(\mreg/_04960_ ), .S(\mreg/_03749_ ), .Z(\mreg/_00315_ ) );
MUX2_X1 \mreg/_09938_ ( .A(\mreg/_04861_ ), .B(\mreg/_04962_ ), .S(\mreg/_03746_ ), .Z(\mreg/_00316_ ) );
MUX2_X1 \mreg/_09939_ ( .A(\mreg/_04862_ ), .B(\mreg/_04963_ ), .S(\mreg/_03746_ ), .Z(\mreg/_00317_ ) );
NAND4_X1 \mreg/_09940_ ( .A1(\mreg/_03691_ ), .A2(\mreg/_03714_ ), .A3(\mreg/_03725_ ), .A4(\mreg/_04937_ ), .ZN(\mreg/_03750_ ) );
NOR2_X1 \mreg/_09941_ ( .A1(\mreg/_03696_ ), .A2(\mreg/_03750_ ), .ZN(\mreg/_03751_ ) );
BUF_X4 \mreg/_09942_ ( .A(\mreg/_03751_ ), .Z(\mreg/_03752_ ) );
MUX2_X1 \mreg/_09943_ ( .A(\mreg/_04870_ ), .B(\mreg/_04939_ ), .S(\mreg/_03752_ ), .Z(\mreg/_00318_ ) );
MUX2_X1 \mreg/_09944_ ( .A(\mreg/_04881_ ), .B(\mreg/_04950_ ), .S(\mreg/_03752_ ), .Z(\mreg/_00319_ ) );
MUX2_X1 \mreg/_09945_ ( .A(\mreg/_04892_ ), .B(\mreg/_04961_ ), .S(\mreg/_03752_ ), .Z(\mreg/_00320_ ) );
MUX2_X1 \mreg/_09946_ ( .A(\mreg/_04895_ ), .B(\mreg/_04964_ ), .S(\mreg/_03752_ ), .Z(\mreg/_00321_ ) );
MUX2_X1 \mreg/_09947_ ( .A(\mreg/_04896_ ), .B(\mreg/_04965_ ), .S(\mreg/_03752_ ), .Z(\mreg/_00322_ ) );
MUX2_X1 \mreg/_09948_ ( .A(\mreg/_04897_ ), .B(\mreg/_04966_ ), .S(\mreg/_03752_ ), .Z(\mreg/_00323_ ) );
MUX2_X1 \mreg/_09949_ ( .A(\mreg/_04898_ ), .B(\mreg/_04967_ ), .S(\mreg/_03752_ ), .Z(\mreg/_00324_ ) );
MUX2_X1 \mreg/_09950_ ( .A(\mreg/_04899_ ), .B(\mreg/_04968_ ), .S(\mreg/_03752_ ), .Z(\mreg/_00325_ ) );
MUX2_X1 \mreg/_09951_ ( .A(\mreg/_04900_ ), .B(\mreg/_04969_ ), .S(\mreg/_03752_ ), .Z(\mreg/_00326_ ) );
MUX2_X1 \mreg/_09952_ ( .A(\mreg/_04901_ ), .B(\mreg/_04970_ ), .S(\mreg/_03752_ ), .Z(\mreg/_00327_ ) );
BUF_X4 \mreg/_09953_ ( .A(\mreg/_03751_ ), .Z(\mreg/_03753_ ) );
MUX2_X1 \mreg/_09954_ ( .A(\mreg/_04871_ ), .B(\mreg/_04940_ ), .S(\mreg/_03753_ ), .Z(\mreg/_00328_ ) );
MUX2_X1 \mreg/_09955_ ( .A(\mreg/_04872_ ), .B(\mreg/_04941_ ), .S(\mreg/_03753_ ), .Z(\mreg/_00329_ ) );
MUX2_X1 \mreg/_09956_ ( .A(\mreg/_04873_ ), .B(\mreg/_04942_ ), .S(\mreg/_03753_ ), .Z(\mreg/_00330_ ) );
MUX2_X1 \mreg/_09957_ ( .A(\mreg/_04874_ ), .B(\mreg/_04943_ ), .S(\mreg/_03753_ ), .Z(\mreg/_00331_ ) );
MUX2_X1 \mreg/_09958_ ( .A(\mreg/_04875_ ), .B(\mreg/_04944_ ), .S(\mreg/_03753_ ), .Z(\mreg/_00332_ ) );
MUX2_X1 \mreg/_09959_ ( .A(\mreg/_04876_ ), .B(\mreg/_04945_ ), .S(\mreg/_03753_ ), .Z(\mreg/_00333_ ) );
MUX2_X1 \mreg/_09960_ ( .A(\mreg/_04877_ ), .B(\mreg/_04946_ ), .S(\mreg/_03753_ ), .Z(\mreg/_00334_ ) );
MUX2_X1 \mreg/_09961_ ( .A(\mreg/_04878_ ), .B(\mreg/_04947_ ), .S(\mreg/_03753_ ), .Z(\mreg/_00335_ ) );
MUX2_X1 \mreg/_09962_ ( .A(\mreg/_04879_ ), .B(\mreg/_04948_ ), .S(\mreg/_03753_ ), .Z(\mreg/_00336_ ) );
MUX2_X1 \mreg/_09963_ ( .A(\mreg/_04880_ ), .B(\mreg/_04949_ ), .S(\mreg/_03753_ ), .Z(\mreg/_00337_ ) );
BUF_X4 \mreg/_09964_ ( .A(\mreg/_03751_ ), .Z(\mreg/_03754_ ) );
MUX2_X1 \mreg/_09965_ ( .A(\mreg/_04882_ ), .B(\mreg/_04951_ ), .S(\mreg/_03754_ ), .Z(\mreg/_00338_ ) );
MUX2_X1 \mreg/_09966_ ( .A(\mreg/_04883_ ), .B(\mreg/_04952_ ), .S(\mreg/_03754_ ), .Z(\mreg/_00339_ ) );
MUX2_X1 \mreg/_09967_ ( .A(\mreg/_04884_ ), .B(\mreg/_04953_ ), .S(\mreg/_03754_ ), .Z(\mreg/_00340_ ) );
MUX2_X1 \mreg/_09968_ ( .A(\mreg/_04885_ ), .B(\mreg/_04954_ ), .S(\mreg/_03754_ ), .Z(\mreg/_00341_ ) );
MUX2_X1 \mreg/_09969_ ( .A(\mreg/_04886_ ), .B(\mreg/_04955_ ), .S(\mreg/_03754_ ), .Z(\mreg/_00342_ ) );
MUX2_X1 \mreg/_09970_ ( .A(\mreg/_04887_ ), .B(\mreg/_04956_ ), .S(\mreg/_03754_ ), .Z(\mreg/_00343_ ) );
MUX2_X1 \mreg/_09971_ ( .A(\mreg/_04888_ ), .B(\mreg/_04957_ ), .S(\mreg/_03754_ ), .Z(\mreg/_00344_ ) );
MUX2_X1 \mreg/_09972_ ( .A(\mreg/_04889_ ), .B(\mreg/_04958_ ), .S(\mreg/_03754_ ), .Z(\mreg/_00345_ ) );
MUX2_X1 \mreg/_09973_ ( .A(\mreg/_04890_ ), .B(\mreg/_04959_ ), .S(\mreg/_03754_ ), .Z(\mreg/_00346_ ) );
MUX2_X1 \mreg/_09974_ ( .A(\mreg/_04891_ ), .B(\mreg/_04960_ ), .S(\mreg/_03754_ ), .Z(\mreg/_00347_ ) );
MUX2_X1 \mreg/_09975_ ( .A(\mreg/_04893_ ), .B(\mreg/_04962_ ), .S(\mreg/_03751_ ), .Z(\mreg/_00348_ ) );
MUX2_X1 \mreg/_09976_ ( .A(\mreg/_04894_ ), .B(\mreg/_04963_ ), .S(\mreg/_03751_ ), .Z(\mreg/_00349_ ) );
NAND2_X1 \mreg/_09977_ ( .A1(\mreg/_03725_ ), .A2(\mreg/_04937_ ), .ZN(\mreg/_03755_ ) );
OR3_X1 \mreg/_09978_ ( .A1(\mreg/_03706_ ), .A2(\mreg/_04938_ ), .A3(\mreg/_03755_ ), .ZN(\mreg/_03756_ ) );
NOR2_X1 \mreg/_09979_ ( .A1(\mreg/_03756_ ), .A2(\mreg/_03709_ ), .ZN(\mreg/_03757_ ) );
BUF_X4 \mreg/_09980_ ( .A(\mreg/_03757_ ), .Z(\mreg/_03758_ ) );
MUX2_X1 \mreg/_09981_ ( .A(\mreg/_04902_ ), .B(\mreg/_04939_ ), .S(\mreg/_03758_ ), .Z(\mreg/_00350_ ) );
MUX2_X1 \mreg/_09982_ ( .A(\mreg/_04913_ ), .B(\mreg/_04950_ ), .S(\mreg/_03758_ ), .Z(\mreg/_00351_ ) );
MUX2_X1 \mreg/_09983_ ( .A(\mreg/_04924_ ), .B(\mreg/_04961_ ), .S(\mreg/_03758_ ), .Z(\mreg/_00352_ ) );
MUX2_X1 \mreg/_09984_ ( .A(\mreg/_04927_ ), .B(\mreg/_04964_ ), .S(\mreg/_03758_ ), .Z(\mreg/_00353_ ) );
MUX2_X1 \mreg/_09985_ ( .A(\mreg/_04928_ ), .B(\mreg/_04965_ ), .S(\mreg/_03758_ ), .Z(\mreg/_00354_ ) );
MUX2_X1 \mreg/_09986_ ( .A(\mreg/_04929_ ), .B(\mreg/_04966_ ), .S(\mreg/_03758_ ), .Z(\mreg/_00355_ ) );
MUX2_X1 \mreg/_09987_ ( .A(\mreg/_04930_ ), .B(\mreg/_04967_ ), .S(\mreg/_03758_ ), .Z(\mreg/_00356_ ) );
MUX2_X1 \mreg/_09988_ ( .A(\mreg/_04931_ ), .B(\mreg/_04968_ ), .S(\mreg/_03758_ ), .Z(\mreg/_00357_ ) );
MUX2_X1 \mreg/_09989_ ( .A(\mreg/_04932_ ), .B(\mreg/_04969_ ), .S(\mreg/_03758_ ), .Z(\mreg/_00358_ ) );
MUX2_X1 \mreg/_09990_ ( .A(\mreg/_04933_ ), .B(\mreg/_04970_ ), .S(\mreg/_03758_ ), .Z(\mreg/_00359_ ) );
BUF_X4 \mreg/_09991_ ( .A(\mreg/_03757_ ), .Z(\mreg/_03759_ ) );
MUX2_X1 \mreg/_09992_ ( .A(\mreg/_04903_ ), .B(\mreg/_04940_ ), .S(\mreg/_03759_ ), .Z(\mreg/_00360_ ) );
MUX2_X1 \mreg/_09993_ ( .A(\mreg/_04904_ ), .B(\mreg/_04941_ ), .S(\mreg/_03759_ ), .Z(\mreg/_00361_ ) );
MUX2_X1 \mreg/_09994_ ( .A(\mreg/_04905_ ), .B(\mreg/_04942_ ), .S(\mreg/_03759_ ), .Z(\mreg/_00362_ ) );
MUX2_X1 \mreg/_09995_ ( .A(\mreg/_04906_ ), .B(\mreg/_04943_ ), .S(\mreg/_03759_ ), .Z(\mreg/_00363_ ) );
MUX2_X1 \mreg/_09996_ ( .A(\mreg/_04907_ ), .B(\mreg/_04944_ ), .S(\mreg/_03759_ ), .Z(\mreg/_00364_ ) );
MUX2_X1 \mreg/_09997_ ( .A(\mreg/_04908_ ), .B(\mreg/_04945_ ), .S(\mreg/_03759_ ), .Z(\mreg/_00365_ ) );
MUX2_X1 \mreg/_09998_ ( .A(\mreg/_04909_ ), .B(\mreg/_04946_ ), .S(\mreg/_03759_ ), .Z(\mreg/_00366_ ) );
MUX2_X1 \mreg/_09999_ ( .A(\mreg/_04910_ ), .B(\mreg/_04947_ ), .S(\mreg/_03759_ ), .Z(\mreg/_00367_ ) );
MUX2_X1 \mreg/_10000_ ( .A(\mreg/_04911_ ), .B(\mreg/_04948_ ), .S(\mreg/_03759_ ), .Z(\mreg/_00368_ ) );
MUX2_X1 \mreg/_10001_ ( .A(\mreg/_04912_ ), .B(\mreg/_04949_ ), .S(\mreg/_03759_ ), .Z(\mreg/_00369_ ) );
BUF_X4 \mreg/_10002_ ( .A(\mreg/_03757_ ), .Z(\mreg/_03760_ ) );
MUX2_X1 \mreg/_10003_ ( .A(\mreg/_04914_ ), .B(\mreg/_04951_ ), .S(\mreg/_03760_ ), .Z(\mreg/_00370_ ) );
MUX2_X1 \mreg/_10004_ ( .A(\mreg/_04915_ ), .B(\mreg/_04952_ ), .S(\mreg/_03760_ ), .Z(\mreg/_00371_ ) );
MUX2_X1 \mreg/_10005_ ( .A(\mreg/_04916_ ), .B(\mreg/_04953_ ), .S(\mreg/_03760_ ), .Z(\mreg/_00372_ ) );
MUX2_X1 \mreg/_10006_ ( .A(\mreg/_04917_ ), .B(\mreg/_04954_ ), .S(\mreg/_03760_ ), .Z(\mreg/_00373_ ) );
MUX2_X1 \mreg/_10007_ ( .A(\mreg/_04918_ ), .B(\mreg/_04955_ ), .S(\mreg/_03760_ ), .Z(\mreg/_00374_ ) );
MUX2_X1 \mreg/_10008_ ( .A(\mreg/_04919_ ), .B(\mreg/_04956_ ), .S(\mreg/_03760_ ), .Z(\mreg/_00375_ ) );
MUX2_X1 \mreg/_10009_ ( .A(\mreg/_04920_ ), .B(\mreg/_04957_ ), .S(\mreg/_03760_ ), .Z(\mreg/_00376_ ) );
MUX2_X1 \mreg/_10010_ ( .A(\mreg/_04921_ ), .B(\mreg/_04958_ ), .S(\mreg/_03760_ ), .Z(\mreg/_00377_ ) );
MUX2_X1 \mreg/_10011_ ( .A(\mreg/_04922_ ), .B(\mreg/_04959_ ), .S(\mreg/_03760_ ), .Z(\mreg/_00378_ ) );
MUX2_X1 \mreg/_10012_ ( .A(\mreg/_04923_ ), .B(\mreg/_04960_ ), .S(\mreg/_03760_ ), .Z(\mreg/_00379_ ) );
MUX2_X1 \mreg/_10013_ ( .A(\mreg/_04925_ ), .B(\mreg/_04962_ ), .S(\mreg/_03757_ ), .Z(\mreg/_00380_ ) );
MUX2_X1 \mreg/_10014_ ( .A(\mreg/_04926_ ), .B(\mreg/_04963_ ), .S(\mreg/_03757_ ), .Z(\mreg/_00381_ ) );
NOR2_X1 \mreg/_10015_ ( .A1(\mreg/_03739_ ), .A2(\mreg/_03755_ ), .ZN(\mreg/_03761_ ) );
NAND2_X1 \mreg/_10016_ ( .A1(\mreg/_03761_ ), .A2(\mreg/_03714_ ), .ZN(\mreg/_03762_ ) );
NOR2_X1 \mreg/_10017_ ( .A1(\mreg/_03762_ ), .A2(\mreg/_03709_ ), .ZN(\mreg/_03763_ ) );
BUF_X4 \mreg/_10018_ ( .A(\mreg/_03763_ ), .Z(\mreg/_03764_ ) );
MUX2_X1 \mreg/_10019_ ( .A(\mreg/_03942_ ), .B(\mreg/_04939_ ), .S(\mreg/_03764_ ), .Z(\mreg/_00382_ ) );
MUX2_X1 \mreg/_10020_ ( .A(\mreg/_03953_ ), .B(\mreg/_04950_ ), .S(\mreg/_03764_ ), .Z(\mreg/_00383_ ) );
MUX2_X1 \mreg/_10021_ ( .A(\mreg/_03964_ ), .B(\mreg/_04961_ ), .S(\mreg/_03764_ ), .Z(\mreg/_00384_ ) );
MUX2_X1 \mreg/_10022_ ( .A(\mreg/_03967_ ), .B(\mreg/_04964_ ), .S(\mreg/_03764_ ), .Z(\mreg/_00385_ ) );
MUX2_X1 \mreg/_10023_ ( .A(\mreg/_03968_ ), .B(\mreg/_04965_ ), .S(\mreg/_03764_ ), .Z(\mreg/_00386_ ) );
MUX2_X1 \mreg/_10024_ ( .A(\mreg/_03969_ ), .B(\mreg/_04966_ ), .S(\mreg/_03764_ ), .Z(\mreg/_00387_ ) );
MUX2_X1 \mreg/_10025_ ( .A(\mreg/_03970_ ), .B(\mreg/_04967_ ), .S(\mreg/_03764_ ), .Z(\mreg/_00388_ ) );
MUX2_X1 \mreg/_10026_ ( .A(\mreg/_03971_ ), .B(\mreg/_04968_ ), .S(\mreg/_03764_ ), .Z(\mreg/_00389_ ) );
MUX2_X1 \mreg/_10027_ ( .A(\mreg/_03972_ ), .B(\mreg/_04969_ ), .S(\mreg/_03764_ ), .Z(\mreg/_00390_ ) );
MUX2_X1 \mreg/_10028_ ( .A(\mreg/_03973_ ), .B(\mreg/_04970_ ), .S(\mreg/_03764_ ), .Z(\mreg/_00391_ ) );
BUF_X4 \mreg/_10029_ ( .A(\mreg/_03763_ ), .Z(\mreg/_03765_ ) );
MUX2_X1 \mreg/_10030_ ( .A(\mreg/_03943_ ), .B(\mreg/_04940_ ), .S(\mreg/_03765_ ), .Z(\mreg/_00392_ ) );
MUX2_X1 \mreg/_10031_ ( .A(\mreg/_03944_ ), .B(\mreg/_04941_ ), .S(\mreg/_03765_ ), .Z(\mreg/_00393_ ) );
MUX2_X1 \mreg/_10032_ ( .A(\mreg/_03945_ ), .B(\mreg/_04942_ ), .S(\mreg/_03765_ ), .Z(\mreg/_00394_ ) );
MUX2_X1 \mreg/_10033_ ( .A(\mreg/_03946_ ), .B(\mreg/_04943_ ), .S(\mreg/_03765_ ), .Z(\mreg/_00395_ ) );
MUX2_X1 \mreg/_10034_ ( .A(\mreg/_03947_ ), .B(\mreg/_04944_ ), .S(\mreg/_03765_ ), .Z(\mreg/_00396_ ) );
MUX2_X1 \mreg/_10035_ ( .A(\mreg/_03948_ ), .B(\mreg/_04945_ ), .S(\mreg/_03765_ ), .Z(\mreg/_00397_ ) );
MUX2_X1 \mreg/_10036_ ( .A(\mreg/_03949_ ), .B(\mreg/_04946_ ), .S(\mreg/_03765_ ), .Z(\mreg/_00398_ ) );
MUX2_X1 \mreg/_10037_ ( .A(\mreg/_03950_ ), .B(\mreg/_04947_ ), .S(\mreg/_03765_ ), .Z(\mreg/_00399_ ) );
MUX2_X1 \mreg/_10038_ ( .A(\mreg/_03951_ ), .B(\mreg/_04948_ ), .S(\mreg/_03765_ ), .Z(\mreg/_00400_ ) );
MUX2_X1 \mreg/_10039_ ( .A(\mreg/_03952_ ), .B(\mreg/_04949_ ), .S(\mreg/_03765_ ), .Z(\mreg/_00401_ ) );
BUF_X4 \mreg/_10040_ ( .A(\mreg/_03763_ ), .Z(\mreg/_03766_ ) );
MUX2_X1 \mreg/_10041_ ( .A(\mreg/_03954_ ), .B(\mreg/_04951_ ), .S(\mreg/_03766_ ), .Z(\mreg/_00402_ ) );
MUX2_X1 \mreg/_10042_ ( .A(\mreg/_03955_ ), .B(\mreg/_04952_ ), .S(\mreg/_03766_ ), .Z(\mreg/_00403_ ) );
MUX2_X1 \mreg/_10043_ ( .A(\mreg/_03956_ ), .B(\mreg/_04953_ ), .S(\mreg/_03766_ ), .Z(\mreg/_00404_ ) );
MUX2_X1 \mreg/_10044_ ( .A(\mreg/_03957_ ), .B(\mreg/_04954_ ), .S(\mreg/_03766_ ), .Z(\mreg/_00405_ ) );
MUX2_X1 \mreg/_10045_ ( .A(\mreg/_03958_ ), .B(\mreg/_04955_ ), .S(\mreg/_03766_ ), .Z(\mreg/_00406_ ) );
MUX2_X1 \mreg/_10046_ ( .A(\mreg/_03959_ ), .B(\mreg/_04956_ ), .S(\mreg/_03766_ ), .Z(\mreg/_00407_ ) );
MUX2_X1 \mreg/_10047_ ( .A(\mreg/_03960_ ), .B(\mreg/_04957_ ), .S(\mreg/_03766_ ), .Z(\mreg/_00408_ ) );
MUX2_X1 \mreg/_10048_ ( .A(\mreg/_03961_ ), .B(\mreg/_04958_ ), .S(\mreg/_03766_ ), .Z(\mreg/_00409_ ) );
MUX2_X1 \mreg/_10049_ ( .A(\mreg/_03962_ ), .B(\mreg/_04959_ ), .S(\mreg/_03766_ ), .Z(\mreg/_00410_ ) );
MUX2_X1 \mreg/_10050_ ( .A(\mreg/_03963_ ), .B(\mreg/_04960_ ), .S(\mreg/_03766_ ), .Z(\mreg/_00411_ ) );
MUX2_X1 \mreg/_10051_ ( .A(\mreg/_03965_ ), .B(\mreg/_04962_ ), .S(\mreg/_03763_ ), .Z(\mreg/_00412_ ) );
MUX2_X1 \mreg/_10052_ ( .A(\mreg/_03966_ ), .B(\mreg/_04963_ ), .S(\mreg/_03763_ ), .Z(\mreg/_00413_ ) );
OR3_X1 \mreg/_10053_ ( .A1(\mreg/_03755_ ), .A2(\mreg/_04938_ ), .A3(\mreg/_03698_ ), .ZN(\mreg/_03767_ ) );
NOR2_X1 \mreg/_10054_ ( .A1(\mreg/_03767_ ), .A2(\mreg/_03709_ ), .ZN(\mreg/_03768_ ) );
BUF_X4 \mreg/_10055_ ( .A(\mreg/_03768_ ), .Z(\mreg/_03769_ ) );
MUX2_X1 \mreg/_10056_ ( .A(\mreg/_03974_ ), .B(\mreg/_04939_ ), .S(\mreg/_03769_ ), .Z(\mreg/_00414_ ) );
MUX2_X1 \mreg/_10057_ ( .A(\mreg/_03985_ ), .B(\mreg/_04950_ ), .S(\mreg/_03769_ ), .Z(\mreg/_00415_ ) );
MUX2_X1 \mreg/_10058_ ( .A(\mreg/_03996_ ), .B(\mreg/_04961_ ), .S(\mreg/_03769_ ), .Z(\mreg/_00416_ ) );
MUX2_X1 \mreg/_10059_ ( .A(\mreg/_03999_ ), .B(\mreg/_04964_ ), .S(\mreg/_03769_ ), .Z(\mreg/_00417_ ) );
MUX2_X1 \mreg/_10060_ ( .A(\mreg/_04000_ ), .B(\mreg/_04965_ ), .S(\mreg/_03769_ ), .Z(\mreg/_00418_ ) );
MUX2_X1 \mreg/_10061_ ( .A(\mreg/_04001_ ), .B(\mreg/_04966_ ), .S(\mreg/_03769_ ), .Z(\mreg/_00419_ ) );
MUX2_X1 \mreg/_10062_ ( .A(\mreg/_04002_ ), .B(\mreg/_04967_ ), .S(\mreg/_03769_ ), .Z(\mreg/_00420_ ) );
MUX2_X1 \mreg/_10063_ ( .A(\mreg/_04003_ ), .B(\mreg/_04968_ ), .S(\mreg/_03769_ ), .Z(\mreg/_00421_ ) );
MUX2_X1 \mreg/_10064_ ( .A(\mreg/_04004_ ), .B(\mreg/_04969_ ), .S(\mreg/_03769_ ), .Z(\mreg/_00422_ ) );
MUX2_X1 \mreg/_10065_ ( .A(\mreg/_04005_ ), .B(\mreg/_04970_ ), .S(\mreg/_03769_ ), .Z(\mreg/_00423_ ) );
BUF_X4 \mreg/_10066_ ( .A(\mreg/_03768_ ), .Z(\mreg/_03770_ ) );
MUX2_X1 \mreg/_10067_ ( .A(\mreg/_03975_ ), .B(\mreg/_04940_ ), .S(\mreg/_03770_ ), .Z(\mreg/_00424_ ) );
MUX2_X1 \mreg/_10068_ ( .A(\mreg/_03976_ ), .B(\mreg/_04941_ ), .S(\mreg/_03770_ ), .Z(\mreg/_00425_ ) );
MUX2_X1 \mreg/_10069_ ( .A(\mreg/_03977_ ), .B(\mreg/_04942_ ), .S(\mreg/_03770_ ), .Z(\mreg/_00426_ ) );
MUX2_X1 \mreg/_10070_ ( .A(\mreg/_03978_ ), .B(\mreg/_04943_ ), .S(\mreg/_03770_ ), .Z(\mreg/_00427_ ) );
MUX2_X1 \mreg/_10071_ ( .A(\mreg/_03979_ ), .B(\mreg/_04944_ ), .S(\mreg/_03770_ ), .Z(\mreg/_00428_ ) );
MUX2_X1 \mreg/_10072_ ( .A(\mreg/_03980_ ), .B(\mreg/_04945_ ), .S(\mreg/_03770_ ), .Z(\mreg/_00429_ ) );
MUX2_X1 \mreg/_10073_ ( .A(\mreg/_03981_ ), .B(\mreg/_04946_ ), .S(\mreg/_03770_ ), .Z(\mreg/_00430_ ) );
MUX2_X1 \mreg/_10074_ ( .A(\mreg/_03982_ ), .B(\mreg/_04947_ ), .S(\mreg/_03770_ ), .Z(\mreg/_00431_ ) );
MUX2_X1 \mreg/_10075_ ( .A(\mreg/_03983_ ), .B(\mreg/_04948_ ), .S(\mreg/_03770_ ), .Z(\mreg/_00432_ ) );
MUX2_X1 \mreg/_10076_ ( .A(\mreg/_03984_ ), .B(\mreg/_04949_ ), .S(\mreg/_03770_ ), .Z(\mreg/_00433_ ) );
BUF_X4 \mreg/_10077_ ( .A(\mreg/_03768_ ), .Z(\mreg/_03771_ ) );
MUX2_X1 \mreg/_10078_ ( .A(\mreg/_03986_ ), .B(\mreg/_04951_ ), .S(\mreg/_03771_ ), .Z(\mreg/_00434_ ) );
MUX2_X1 \mreg/_10079_ ( .A(\mreg/_03987_ ), .B(\mreg/_04952_ ), .S(\mreg/_03771_ ), .Z(\mreg/_00435_ ) );
MUX2_X1 \mreg/_10080_ ( .A(\mreg/_03988_ ), .B(\mreg/_04953_ ), .S(\mreg/_03771_ ), .Z(\mreg/_00436_ ) );
MUX2_X1 \mreg/_10081_ ( .A(\mreg/_03989_ ), .B(\mreg/_04954_ ), .S(\mreg/_03771_ ), .Z(\mreg/_00437_ ) );
MUX2_X1 \mreg/_10082_ ( .A(\mreg/_03990_ ), .B(\mreg/_04955_ ), .S(\mreg/_03771_ ), .Z(\mreg/_00438_ ) );
MUX2_X1 \mreg/_10083_ ( .A(\mreg/_03991_ ), .B(\mreg/_04956_ ), .S(\mreg/_03771_ ), .Z(\mreg/_00439_ ) );
MUX2_X1 \mreg/_10084_ ( .A(\mreg/_03992_ ), .B(\mreg/_04957_ ), .S(\mreg/_03771_ ), .Z(\mreg/_00440_ ) );
MUX2_X1 \mreg/_10085_ ( .A(\mreg/_03993_ ), .B(\mreg/_04958_ ), .S(\mreg/_03771_ ), .Z(\mreg/_00441_ ) );
MUX2_X1 \mreg/_10086_ ( .A(\mreg/_03994_ ), .B(\mreg/_04959_ ), .S(\mreg/_03771_ ), .Z(\mreg/_00442_ ) );
MUX2_X1 \mreg/_10087_ ( .A(\mreg/_03995_ ), .B(\mreg/_04960_ ), .S(\mreg/_03771_ ), .Z(\mreg/_00443_ ) );
MUX2_X1 \mreg/_10088_ ( .A(\mreg/_03997_ ), .B(\mreg/_04962_ ), .S(\mreg/_03768_ ), .Z(\mreg/_00444_ ) );
MUX2_X1 \mreg/_10089_ ( .A(\mreg/_03998_ ), .B(\mreg/_04963_ ), .S(\mreg/_03768_ ), .Z(\mreg/_00445_ ) );
NAND4_X1 \mreg/_10090_ ( .A1(\mreg/_03691_ ), .A2(\mreg/_03714_ ), .A3(\mreg/_04936_ ), .A4(\mreg/_04937_ ), .ZN(\mreg/_03772_ ) );
NOR2_X1 \mreg/_10091_ ( .A1(\mreg/_03696_ ), .A2(\mreg/_03772_ ), .ZN(\mreg/_03773_ ) );
BUF_X4 \mreg/_10092_ ( .A(\mreg/_03773_ ), .Z(\mreg/_03774_ ) );
MUX2_X1 \mreg/_10093_ ( .A(\mreg/_04006_ ), .B(\mreg/_04939_ ), .S(\mreg/_03774_ ), .Z(\mreg/_00446_ ) );
MUX2_X1 \mreg/_10094_ ( .A(\mreg/_04017_ ), .B(\mreg/_04950_ ), .S(\mreg/_03774_ ), .Z(\mreg/_00447_ ) );
MUX2_X1 \mreg/_10095_ ( .A(\mreg/_04028_ ), .B(\mreg/_04961_ ), .S(\mreg/_03774_ ), .Z(\mreg/_00448_ ) );
MUX2_X1 \mreg/_10096_ ( .A(\mreg/_04031_ ), .B(\mreg/_04964_ ), .S(\mreg/_03774_ ), .Z(\mreg/_00449_ ) );
MUX2_X1 \mreg/_10097_ ( .A(\mreg/_04032_ ), .B(\mreg/_04965_ ), .S(\mreg/_03774_ ), .Z(\mreg/_00450_ ) );
MUX2_X1 \mreg/_10098_ ( .A(\mreg/_04033_ ), .B(\mreg/_04966_ ), .S(\mreg/_03774_ ), .Z(\mreg/_00451_ ) );
MUX2_X1 \mreg/_10099_ ( .A(\mreg/_04034_ ), .B(\mreg/_04967_ ), .S(\mreg/_03774_ ), .Z(\mreg/_00452_ ) );
MUX2_X1 \mreg/_10100_ ( .A(\mreg/_04035_ ), .B(\mreg/_04968_ ), .S(\mreg/_03774_ ), .Z(\mreg/_00453_ ) );
MUX2_X1 \mreg/_10101_ ( .A(\mreg/_04036_ ), .B(\mreg/_04969_ ), .S(\mreg/_03774_ ), .Z(\mreg/_00454_ ) );
MUX2_X1 \mreg/_10102_ ( .A(\mreg/_04037_ ), .B(\mreg/_04970_ ), .S(\mreg/_03774_ ), .Z(\mreg/_00455_ ) );
BUF_X4 \mreg/_10103_ ( .A(\mreg/_03773_ ), .Z(\mreg/_03775_ ) );
MUX2_X1 \mreg/_10104_ ( .A(\mreg/_04007_ ), .B(\mreg/_04940_ ), .S(\mreg/_03775_ ), .Z(\mreg/_00456_ ) );
MUX2_X1 \mreg/_10105_ ( .A(\mreg/_04008_ ), .B(\mreg/_04941_ ), .S(\mreg/_03775_ ), .Z(\mreg/_00457_ ) );
MUX2_X1 \mreg/_10106_ ( .A(\mreg/_04009_ ), .B(\mreg/_04942_ ), .S(\mreg/_03775_ ), .Z(\mreg/_00458_ ) );
MUX2_X1 \mreg/_10107_ ( .A(\mreg/_04010_ ), .B(\mreg/_04943_ ), .S(\mreg/_03775_ ), .Z(\mreg/_00459_ ) );
MUX2_X1 \mreg/_10108_ ( .A(\mreg/_04011_ ), .B(\mreg/_04944_ ), .S(\mreg/_03775_ ), .Z(\mreg/_00460_ ) );
MUX2_X1 \mreg/_10109_ ( .A(\mreg/_04012_ ), .B(\mreg/_04945_ ), .S(\mreg/_03775_ ), .Z(\mreg/_00461_ ) );
MUX2_X1 \mreg/_10110_ ( .A(\mreg/_04013_ ), .B(\mreg/_04946_ ), .S(\mreg/_03775_ ), .Z(\mreg/_00462_ ) );
MUX2_X1 \mreg/_10111_ ( .A(\mreg/_04014_ ), .B(\mreg/_04947_ ), .S(\mreg/_03775_ ), .Z(\mreg/_00463_ ) );
MUX2_X1 \mreg/_10112_ ( .A(\mreg/_04015_ ), .B(\mreg/_04948_ ), .S(\mreg/_03775_ ), .Z(\mreg/_00464_ ) );
MUX2_X1 \mreg/_10113_ ( .A(\mreg/_04016_ ), .B(\mreg/_04949_ ), .S(\mreg/_03775_ ), .Z(\mreg/_00465_ ) );
BUF_X4 \mreg/_10114_ ( .A(\mreg/_03773_ ), .Z(\mreg/_03776_ ) );
MUX2_X1 \mreg/_10115_ ( .A(\mreg/_04018_ ), .B(\mreg/_04951_ ), .S(\mreg/_03776_ ), .Z(\mreg/_00466_ ) );
MUX2_X1 \mreg/_10116_ ( .A(\mreg/_04019_ ), .B(\mreg/_04952_ ), .S(\mreg/_03776_ ), .Z(\mreg/_00467_ ) );
MUX2_X1 \mreg/_10117_ ( .A(\mreg/_04020_ ), .B(\mreg/_04953_ ), .S(\mreg/_03776_ ), .Z(\mreg/_00468_ ) );
MUX2_X1 \mreg/_10118_ ( .A(\mreg/_04021_ ), .B(\mreg/_04954_ ), .S(\mreg/_03776_ ), .Z(\mreg/_00469_ ) );
MUX2_X1 \mreg/_10119_ ( .A(\mreg/_04022_ ), .B(\mreg/_04955_ ), .S(\mreg/_03776_ ), .Z(\mreg/_00470_ ) );
MUX2_X1 \mreg/_10120_ ( .A(\mreg/_04023_ ), .B(\mreg/_04956_ ), .S(\mreg/_03776_ ), .Z(\mreg/_00471_ ) );
MUX2_X1 \mreg/_10121_ ( .A(\mreg/_04024_ ), .B(\mreg/_04957_ ), .S(\mreg/_03776_ ), .Z(\mreg/_00472_ ) );
MUX2_X1 \mreg/_10122_ ( .A(\mreg/_04025_ ), .B(\mreg/_04958_ ), .S(\mreg/_03776_ ), .Z(\mreg/_00473_ ) );
MUX2_X1 \mreg/_10123_ ( .A(\mreg/_04026_ ), .B(\mreg/_04959_ ), .S(\mreg/_03776_ ), .Z(\mreg/_00474_ ) );
MUX2_X1 \mreg/_10124_ ( .A(\mreg/_04027_ ), .B(\mreg/_04960_ ), .S(\mreg/_03776_ ), .Z(\mreg/_00475_ ) );
MUX2_X1 \mreg/_10125_ ( .A(\mreg/_04029_ ), .B(\mreg/_04962_ ), .S(\mreg/_03773_ ), .Z(\mreg/_00476_ ) );
MUX2_X1 \mreg/_10126_ ( .A(\mreg/_04030_ ), .B(\mreg/_04963_ ), .S(\mreg/_03773_ ), .Z(\mreg/_00477_ ) );
OR4_X1 \mreg/_10127_ ( .A1(\mreg/_04938_ ), .A2(\mreg/_03697_ ), .A3(\mreg/_03705_ ), .A4(\mreg/_04935_ ), .ZN(\mreg/_03777_ ) );
NOR2_X1 \mreg/_10128_ ( .A1(\mreg/_03777_ ), .A2(\mreg/_03709_ ), .ZN(\mreg/_03778_ ) );
BUF_X4 \mreg/_10129_ ( .A(\mreg/_03778_ ), .Z(\mreg/_03779_ ) );
MUX2_X1 \mreg/_10130_ ( .A(\mreg/_04038_ ), .B(\mreg/_04939_ ), .S(\mreg/_03779_ ), .Z(\mreg/_00478_ ) );
MUX2_X1 \mreg/_10131_ ( .A(\mreg/_04049_ ), .B(\mreg/_04950_ ), .S(\mreg/_03779_ ), .Z(\mreg/_00479_ ) );
MUX2_X1 \mreg/_10132_ ( .A(\mreg/_04060_ ), .B(\mreg/_04961_ ), .S(\mreg/_03779_ ), .Z(\mreg/_00480_ ) );
MUX2_X1 \mreg/_10133_ ( .A(\mreg/_04063_ ), .B(\mreg/_04964_ ), .S(\mreg/_03779_ ), .Z(\mreg/_00481_ ) );
MUX2_X1 \mreg/_10134_ ( .A(\mreg/_04064_ ), .B(\mreg/_04965_ ), .S(\mreg/_03779_ ), .Z(\mreg/_00482_ ) );
MUX2_X1 \mreg/_10135_ ( .A(\mreg/_04065_ ), .B(\mreg/_04966_ ), .S(\mreg/_03779_ ), .Z(\mreg/_00483_ ) );
MUX2_X1 \mreg/_10136_ ( .A(\mreg/_04066_ ), .B(\mreg/_04967_ ), .S(\mreg/_03779_ ), .Z(\mreg/_00484_ ) );
MUX2_X1 \mreg/_10137_ ( .A(\mreg/_04067_ ), .B(\mreg/_04968_ ), .S(\mreg/_03779_ ), .Z(\mreg/_00485_ ) );
MUX2_X1 \mreg/_10138_ ( .A(\mreg/_04068_ ), .B(\mreg/_04969_ ), .S(\mreg/_03779_ ), .Z(\mreg/_00486_ ) );
MUX2_X1 \mreg/_10139_ ( .A(\mreg/_04069_ ), .B(\mreg/_04970_ ), .S(\mreg/_03779_ ), .Z(\mreg/_00487_ ) );
BUF_X4 \mreg/_10140_ ( .A(\mreg/_03778_ ), .Z(\mreg/_03780_ ) );
MUX2_X1 \mreg/_10141_ ( .A(\mreg/_04039_ ), .B(\mreg/_04940_ ), .S(\mreg/_03780_ ), .Z(\mreg/_00488_ ) );
MUX2_X1 \mreg/_10142_ ( .A(\mreg/_04040_ ), .B(\mreg/_04941_ ), .S(\mreg/_03780_ ), .Z(\mreg/_00489_ ) );
MUX2_X1 \mreg/_10143_ ( .A(\mreg/_04041_ ), .B(\mreg/_04942_ ), .S(\mreg/_03780_ ), .Z(\mreg/_00490_ ) );
MUX2_X1 \mreg/_10144_ ( .A(\mreg/_04042_ ), .B(\mreg/_04943_ ), .S(\mreg/_03780_ ), .Z(\mreg/_00491_ ) );
MUX2_X1 \mreg/_10145_ ( .A(\mreg/_04043_ ), .B(\mreg/_04944_ ), .S(\mreg/_03780_ ), .Z(\mreg/_00492_ ) );
MUX2_X1 \mreg/_10146_ ( .A(\mreg/_04044_ ), .B(\mreg/_04945_ ), .S(\mreg/_03780_ ), .Z(\mreg/_00493_ ) );
MUX2_X1 \mreg/_10147_ ( .A(\mreg/_04045_ ), .B(\mreg/_04946_ ), .S(\mreg/_03780_ ), .Z(\mreg/_00494_ ) );
MUX2_X1 \mreg/_10148_ ( .A(\mreg/_04046_ ), .B(\mreg/_04947_ ), .S(\mreg/_03780_ ), .Z(\mreg/_00495_ ) );
MUX2_X1 \mreg/_10149_ ( .A(\mreg/_04047_ ), .B(\mreg/_04948_ ), .S(\mreg/_03780_ ), .Z(\mreg/_00496_ ) );
MUX2_X1 \mreg/_10150_ ( .A(\mreg/_04048_ ), .B(\mreg/_04949_ ), .S(\mreg/_03780_ ), .Z(\mreg/_00497_ ) );
BUF_X4 \mreg/_10151_ ( .A(\mreg/_03778_ ), .Z(\mreg/_03781_ ) );
MUX2_X1 \mreg/_10152_ ( .A(\mreg/_04050_ ), .B(\mreg/_04951_ ), .S(\mreg/_03781_ ), .Z(\mreg/_00498_ ) );
MUX2_X1 \mreg/_10153_ ( .A(\mreg/_04051_ ), .B(\mreg/_04952_ ), .S(\mreg/_03781_ ), .Z(\mreg/_00499_ ) );
MUX2_X1 \mreg/_10154_ ( .A(\mreg/_04052_ ), .B(\mreg/_04953_ ), .S(\mreg/_03781_ ), .Z(\mreg/_00500_ ) );
MUX2_X1 \mreg/_10155_ ( .A(\mreg/_04053_ ), .B(\mreg/_04954_ ), .S(\mreg/_03781_ ), .Z(\mreg/_00501_ ) );
MUX2_X1 \mreg/_10156_ ( .A(\mreg/_04054_ ), .B(\mreg/_04955_ ), .S(\mreg/_03781_ ), .Z(\mreg/_00502_ ) );
MUX2_X1 \mreg/_10157_ ( .A(\mreg/_04055_ ), .B(\mreg/_04956_ ), .S(\mreg/_03781_ ), .Z(\mreg/_00503_ ) );
MUX2_X1 \mreg/_10158_ ( .A(\mreg/_04056_ ), .B(\mreg/_04957_ ), .S(\mreg/_03781_ ), .Z(\mreg/_00504_ ) );
MUX2_X1 \mreg/_10159_ ( .A(\mreg/_04057_ ), .B(\mreg/_04958_ ), .S(\mreg/_03781_ ), .Z(\mreg/_00505_ ) );
MUX2_X1 \mreg/_10160_ ( .A(\mreg/_04058_ ), .B(\mreg/_04959_ ), .S(\mreg/_03781_ ), .Z(\mreg/_00506_ ) );
MUX2_X1 \mreg/_10161_ ( .A(\mreg/_04059_ ), .B(\mreg/_04960_ ), .S(\mreg/_03781_ ), .Z(\mreg/_00507_ ) );
MUX2_X1 \mreg/_10162_ ( .A(\mreg/_04061_ ), .B(\mreg/_04962_ ), .S(\mreg/_03778_ ), .Z(\mreg/_00508_ ) );
MUX2_X1 \mreg/_10163_ ( .A(\mreg/_04062_ ), .B(\mreg/_04963_ ), .S(\mreg/_03778_ ), .Z(\mreg/_00509_ ) );
OR3_X1 \mreg/_10164_ ( .A1(\mreg/_03739_ ), .A2(\mreg/_04938_ ), .A3(\mreg/_03697_ ), .ZN(\mreg/_03782_ ) );
BUF_X4 \mreg/_10165_ ( .A(\mreg/_03695_ ), .Z(\mreg/_03783_ ) );
NOR2_X1 \mreg/_10166_ ( .A1(\mreg/_03782_ ), .A2(\mreg/_03783_ ), .ZN(\mreg/_03784_ ) );
BUF_X4 \mreg/_10167_ ( .A(\mreg/_03784_ ), .Z(\mreg/_03785_ ) );
MUX2_X1 \mreg/_10168_ ( .A(\mreg/_04070_ ), .B(\mreg/_04939_ ), .S(\mreg/_03785_ ), .Z(\mreg/_00510_ ) );
MUX2_X1 \mreg/_10169_ ( .A(\mreg/_04081_ ), .B(\mreg/_04950_ ), .S(\mreg/_03785_ ), .Z(\mreg/_00511_ ) );
MUX2_X1 \mreg/_10170_ ( .A(\mreg/_04092_ ), .B(\mreg/_04961_ ), .S(\mreg/_03785_ ), .Z(\mreg/_00512_ ) );
MUX2_X1 \mreg/_10171_ ( .A(\mreg/_04095_ ), .B(\mreg/_04964_ ), .S(\mreg/_03785_ ), .Z(\mreg/_00513_ ) );
MUX2_X1 \mreg/_10172_ ( .A(\mreg/_04096_ ), .B(\mreg/_04965_ ), .S(\mreg/_03785_ ), .Z(\mreg/_00514_ ) );
MUX2_X1 \mreg/_10173_ ( .A(\mreg/_04097_ ), .B(\mreg/_04966_ ), .S(\mreg/_03785_ ), .Z(\mreg/_00515_ ) );
MUX2_X1 \mreg/_10174_ ( .A(\mreg/_04098_ ), .B(\mreg/_04967_ ), .S(\mreg/_03785_ ), .Z(\mreg/_00516_ ) );
MUX2_X1 \mreg/_10175_ ( .A(\mreg/_04099_ ), .B(\mreg/_04968_ ), .S(\mreg/_03785_ ), .Z(\mreg/_00517_ ) );
MUX2_X1 \mreg/_10176_ ( .A(\mreg/_04100_ ), .B(\mreg/_04969_ ), .S(\mreg/_03785_ ), .Z(\mreg/_00518_ ) );
MUX2_X1 \mreg/_10177_ ( .A(\mreg/_04101_ ), .B(\mreg/_04970_ ), .S(\mreg/_03785_ ), .Z(\mreg/_00519_ ) );
BUF_X4 \mreg/_10178_ ( .A(\mreg/_03784_ ), .Z(\mreg/_03786_ ) );
MUX2_X1 \mreg/_10179_ ( .A(\mreg/_04071_ ), .B(\mreg/_04940_ ), .S(\mreg/_03786_ ), .Z(\mreg/_00520_ ) );
MUX2_X1 \mreg/_10180_ ( .A(\mreg/_04072_ ), .B(\mreg/_04941_ ), .S(\mreg/_03786_ ), .Z(\mreg/_00521_ ) );
MUX2_X1 \mreg/_10181_ ( .A(\mreg/_04073_ ), .B(\mreg/_04942_ ), .S(\mreg/_03786_ ), .Z(\mreg/_00522_ ) );
MUX2_X1 \mreg/_10182_ ( .A(\mreg/_04074_ ), .B(\mreg/_04943_ ), .S(\mreg/_03786_ ), .Z(\mreg/_00523_ ) );
MUX2_X1 \mreg/_10183_ ( .A(\mreg/_04075_ ), .B(\mreg/_04944_ ), .S(\mreg/_03786_ ), .Z(\mreg/_00524_ ) );
MUX2_X1 \mreg/_10184_ ( .A(\mreg/_04076_ ), .B(\mreg/_04945_ ), .S(\mreg/_03786_ ), .Z(\mreg/_00525_ ) );
MUX2_X1 \mreg/_10185_ ( .A(\mreg/_04077_ ), .B(\mreg/_04946_ ), .S(\mreg/_03786_ ), .Z(\mreg/_00526_ ) );
MUX2_X1 \mreg/_10186_ ( .A(\mreg/_04078_ ), .B(\mreg/_04947_ ), .S(\mreg/_03786_ ), .Z(\mreg/_00527_ ) );
MUX2_X1 \mreg/_10187_ ( .A(\mreg/_04079_ ), .B(\mreg/_04948_ ), .S(\mreg/_03786_ ), .Z(\mreg/_00528_ ) );
MUX2_X1 \mreg/_10188_ ( .A(\mreg/_04080_ ), .B(\mreg/_04949_ ), .S(\mreg/_03786_ ), .Z(\mreg/_00529_ ) );
BUF_X4 \mreg/_10189_ ( .A(\mreg/_03784_ ), .Z(\mreg/_03787_ ) );
MUX2_X1 \mreg/_10190_ ( .A(\mreg/_04082_ ), .B(\mreg/_04951_ ), .S(\mreg/_03787_ ), .Z(\mreg/_00530_ ) );
MUX2_X1 \mreg/_10191_ ( .A(\mreg/_04083_ ), .B(\mreg/_04952_ ), .S(\mreg/_03787_ ), .Z(\mreg/_00531_ ) );
MUX2_X1 \mreg/_10192_ ( .A(\mreg/_04084_ ), .B(\mreg/_04953_ ), .S(\mreg/_03787_ ), .Z(\mreg/_00532_ ) );
MUX2_X1 \mreg/_10193_ ( .A(\mreg/_04085_ ), .B(\mreg/_04954_ ), .S(\mreg/_03787_ ), .Z(\mreg/_00533_ ) );
MUX2_X1 \mreg/_10194_ ( .A(\mreg/_04086_ ), .B(\mreg/_04955_ ), .S(\mreg/_03787_ ), .Z(\mreg/_00534_ ) );
MUX2_X1 \mreg/_10195_ ( .A(\mreg/_04087_ ), .B(\mreg/_04956_ ), .S(\mreg/_03787_ ), .Z(\mreg/_00535_ ) );
MUX2_X1 \mreg/_10196_ ( .A(\mreg/_04088_ ), .B(\mreg/_04957_ ), .S(\mreg/_03787_ ), .Z(\mreg/_00536_ ) );
MUX2_X1 \mreg/_10197_ ( .A(\mreg/_04089_ ), .B(\mreg/_04958_ ), .S(\mreg/_03787_ ), .Z(\mreg/_00537_ ) );
MUX2_X1 \mreg/_10198_ ( .A(\mreg/_04090_ ), .B(\mreg/_04959_ ), .S(\mreg/_03787_ ), .Z(\mreg/_00538_ ) );
MUX2_X1 \mreg/_10199_ ( .A(\mreg/_04091_ ), .B(\mreg/_04960_ ), .S(\mreg/_03787_ ), .Z(\mreg/_00539_ ) );
MUX2_X1 \mreg/_10200_ ( .A(\mreg/_04093_ ), .B(\mreg/_04962_ ), .S(\mreg/_03784_ ), .Z(\mreg/_00540_ ) );
MUX2_X1 \mreg/_10201_ ( .A(\mreg/_04094_ ), .B(\mreg/_04963_ ), .S(\mreg/_03784_ ), .Z(\mreg/_00541_ ) );
NAND2_X1 \mreg/_10202_ ( .A1(\mreg/_03699_ ), .A2(\mreg/_03714_ ), .ZN(\mreg/_03788_ ) );
NOR2_X1 \mreg/_10203_ ( .A1(\mreg/_03696_ ), .A2(\mreg/_03788_ ), .ZN(\mreg/_03789_ ) );
BUF_X4 \mreg/_10204_ ( .A(\mreg/_03789_ ), .Z(\mreg/_03790_ ) );
MUX2_X1 \mreg/_10205_ ( .A(\mreg/_04102_ ), .B(\mreg/_04939_ ), .S(\mreg/_03790_ ), .Z(\mreg/_00542_ ) );
MUX2_X1 \mreg/_10206_ ( .A(\mreg/_04113_ ), .B(\mreg/_04950_ ), .S(\mreg/_03790_ ), .Z(\mreg/_00543_ ) );
MUX2_X1 \mreg/_10207_ ( .A(\mreg/_04124_ ), .B(\mreg/_04961_ ), .S(\mreg/_03790_ ), .Z(\mreg/_00544_ ) );
MUX2_X1 \mreg/_10208_ ( .A(\mreg/_04127_ ), .B(\mreg/_04964_ ), .S(\mreg/_03790_ ), .Z(\mreg/_00545_ ) );
MUX2_X1 \mreg/_10209_ ( .A(\mreg/_04128_ ), .B(\mreg/_04965_ ), .S(\mreg/_03790_ ), .Z(\mreg/_00546_ ) );
MUX2_X1 \mreg/_10210_ ( .A(\mreg/_04129_ ), .B(\mreg/_04966_ ), .S(\mreg/_03790_ ), .Z(\mreg/_00547_ ) );
MUX2_X1 \mreg/_10211_ ( .A(\mreg/_04130_ ), .B(\mreg/_04967_ ), .S(\mreg/_03790_ ), .Z(\mreg/_00548_ ) );
MUX2_X1 \mreg/_10212_ ( .A(\mreg/_04131_ ), .B(\mreg/_04968_ ), .S(\mreg/_03790_ ), .Z(\mreg/_00549_ ) );
MUX2_X1 \mreg/_10213_ ( .A(\mreg/_04132_ ), .B(\mreg/_04969_ ), .S(\mreg/_03790_ ), .Z(\mreg/_00550_ ) );
MUX2_X1 \mreg/_10214_ ( .A(\mreg/_04133_ ), .B(\mreg/_04970_ ), .S(\mreg/_03790_ ), .Z(\mreg/_00551_ ) );
BUF_X4 \mreg/_10215_ ( .A(\mreg/_03789_ ), .Z(\mreg/_03791_ ) );
MUX2_X1 \mreg/_10216_ ( .A(\mreg/_04103_ ), .B(\mreg/_04940_ ), .S(\mreg/_03791_ ), .Z(\mreg/_00552_ ) );
MUX2_X1 \mreg/_10217_ ( .A(\mreg/_04104_ ), .B(\mreg/_04941_ ), .S(\mreg/_03791_ ), .Z(\mreg/_00553_ ) );
MUX2_X1 \mreg/_10218_ ( .A(\mreg/_04105_ ), .B(\mreg/_04942_ ), .S(\mreg/_03791_ ), .Z(\mreg/_00554_ ) );
MUX2_X1 \mreg/_10219_ ( .A(\mreg/_04106_ ), .B(\mreg/_04943_ ), .S(\mreg/_03791_ ), .Z(\mreg/_00555_ ) );
MUX2_X1 \mreg/_10220_ ( .A(\mreg/_04107_ ), .B(\mreg/_04944_ ), .S(\mreg/_03791_ ), .Z(\mreg/_00556_ ) );
MUX2_X1 \mreg/_10221_ ( .A(\mreg/_04108_ ), .B(\mreg/_04945_ ), .S(\mreg/_03791_ ), .Z(\mreg/_00557_ ) );
MUX2_X1 \mreg/_10222_ ( .A(\mreg/_04109_ ), .B(\mreg/_04946_ ), .S(\mreg/_03791_ ), .Z(\mreg/_00558_ ) );
MUX2_X1 \mreg/_10223_ ( .A(\mreg/_04110_ ), .B(\mreg/_04947_ ), .S(\mreg/_03791_ ), .Z(\mreg/_00559_ ) );
MUX2_X1 \mreg/_10224_ ( .A(\mreg/_04111_ ), .B(\mreg/_04948_ ), .S(\mreg/_03791_ ), .Z(\mreg/_00560_ ) );
MUX2_X1 \mreg/_10225_ ( .A(\mreg/_04112_ ), .B(\mreg/_04949_ ), .S(\mreg/_03791_ ), .Z(\mreg/_00561_ ) );
BUF_X4 \mreg/_10226_ ( .A(\mreg/_03789_ ), .Z(\mreg/_03792_ ) );
MUX2_X1 \mreg/_10227_ ( .A(\mreg/_04114_ ), .B(\mreg/_04951_ ), .S(\mreg/_03792_ ), .Z(\mreg/_00562_ ) );
MUX2_X1 \mreg/_10228_ ( .A(\mreg/_04115_ ), .B(\mreg/_04952_ ), .S(\mreg/_03792_ ), .Z(\mreg/_00563_ ) );
MUX2_X1 \mreg/_10229_ ( .A(\mreg/_04116_ ), .B(\mreg/_04953_ ), .S(\mreg/_03792_ ), .Z(\mreg/_00564_ ) );
MUX2_X1 \mreg/_10230_ ( .A(\mreg/_04117_ ), .B(\mreg/_04954_ ), .S(\mreg/_03792_ ), .Z(\mreg/_00565_ ) );
MUX2_X1 \mreg/_10231_ ( .A(\mreg/_04118_ ), .B(\mreg/_04955_ ), .S(\mreg/_03792_ ), .Z(\mreg/_00566_ ) );
MUX2_X1 \mreg/_10232_ ( .A(\mreg/_04119_ ), .B(\mreg/_04956_ ), .S(\mreg/_03792_ ), .Z(\mreg/_00567_ ) );
MUX2_X1 \mreg/_10233_ ( .A(\mreg/_04120_ ), .B(\mreg/_04957_ ), .S(\mreg/_03792_ ), .Z(\mreg/_00568_ ) );
MUX2_X1 \mreg/_10234_ ( .A(\mreg/_04121_ ), .B(\mreg/_04958_ ), .S(\mreg/_03792_ ), .Z(\mreg/_00569_ ) );
MUX2_X1 \mreg/_10235_ ( .A(\mreg/_04122_ ), .B(\mreg/_04959_ ), .S(\mreg/_03792_ ), .Z(\mreg/_00570_ ) );
MUX2_X1 \mreg/_10236_ ( .A(\mreg/_04123_ ), .B(\mreg/_04960_ ), .S(\mreg/_03792_ ), .Z(\mreg/_00571_ ) );
MUX2_X1 \mreg/_10237_ ( .A(\mreg/_04125_ ), .B(\mreg/_04962_ ), .S(\mreg/_03789_ ), .Z(\mreg/_00572_ ) );
MUX2_X1 \mreg/_10238_ ( .A(\mreg/_04126_ ), .B(\mreg/_04963_ ), .S(\mreg/_03789_ ), .Z(\mreg/_00573_ ) );
NAND3_X1 \mreg/_10239_ ( .A1(\mreg/_03690_ ), .A2(\mreg/_03691_ ), .A3(\mreg/_04938_ ), .ZN(\mreg/_03793_ ) );
NOR2_X1 \mreg/_10240_ ( .A1(\mreg/_03696_ ), .A2(\mreg/_03793_ ), .ZN(\mreg/_03794_ ) );
BUF_X4 \mreg/_10241_ ( .A(\mreg/_03794_ ), .Z(\mreg/_03795_ ) );
MUX2_X1 \mreg/_10242_ ( .A(\mreg/_04134_ ), .B(\mreg/_04939_ ), .S(\mreg/_03795_ ), .Z(\mreg/_00574_ ) );
MUX2_X1 \mreg/_10243_ ( .A(\mreg/_04145_ ), .B(\mreg/_04950_ ), .S(\mreg/_03795_ ), .Z(\mreg/_00575_ ) );
MUX2_X1 \mreg/_10244_ ( .A(\mreg/_04156_ ), .B(\mreg/_04961_ ), .S(\mreg/_03795_ ), .Z(\mreg/_00576_ ) );
MUX2_X1 \mreg/_10245_ ( .A(\mreg/_04159_ ), .B(\mreg/_04964_ ), .S(\mreg/_03795_ ), .Z(\mreg/_00577_ ) );
MUX2_X1 \mreg/_10246_ ( .A(\mreg/_04160_ ), .B(\mreg/_04965_ ), .S(\mreg/_03795_ ), .Z(\mreg/_00578_ ) );
MUX2_X1 \mreg/_10247_ ( .A(\mreg/_04161_ ), .B(\mreg/_04966_ ), .S(\mreg/_03795_ ), .Z(\mreg/_00579_ ) );
MUX2_X1 \mreg/_10248_ ( .A(\mreg/_04162_ ), .B(\mreg/_04967_ ), .S(\mreg/_03795_ ), .Z(\mreg/_00580_ ) );
MUX2_X1 \mreg/_10249_ ( .A(\mreg/_04163_ ), .B(\mreg/_04968_ ), .S(\mreg/_03795_ ), .Z(\mreg/_00581_ ) );
MUX2_X1 \mreg/_10250_ ( .A(\mreg/_04164_ ), .B(\mreg/_04969_ ), .S(\mreg/_03795_ ), .Z(\mreg/_00582_ ) );
MUX2_X1 \mreg/_10251_ ( .A(\mreg/_04165_ ), .B(\mreg/_04970_ ), .S(\mreg/_03795_ ), .Z(\mreg/_00583_ ) );
BUF_X4 \mreg/_10252_ ( .A(\mreg/_03794_ ), .Z(\mreg/_03796_ ) );
MUX2_X1 \mreg/_10253_ ( .A(\mreg/_04135_ ), .B(\mreg/_04940_ ), .S(\mreg/_03796_ ), .Z(\mreg/_00584_ ) );
MUX2_X1 \mreg/_10254_ ( .A(\mreg/_04136_ ), .B(\mreg/_04941_ ), .S(\mreg/_03796_ ), .Z(\mreg/_00585_ ) );
MUX2_X1 \mreg/_10255_ ( .A(\mreg/_04137_ ), .B(\mreg/_04942_ ), .S(\mreg/_03796_ ), .Z(\mreg/_00586_ ) );
MUX2_X1 \mreg/_10256_ ( .A(\mreg/_04138_ ), .B(\mreg/_04943_ ), .S(\mreg/_03796_ ), .Z(\mreg/_00587_ ) );
MUX2_X1 \mreg/_10257_ ( .A(\mreg/_04139_ ), .B(\mreg/_04944_ ), .S(\mreg/_03796_ ), .Z(\mreg/_00588_ ) );
MUX2_X1 \mreg/_10258_ ( .A(\mreg/_04140_ ), .B(\mreg/_04945_ ), .S(\mreg/_03796_ ), .Z(\mreg/_00589_ ) );
MUX2_X1 \mreg/_10259_ ( .A(\mreg/_04141_ ), .B(\mreg/_04946_ ), .S(\mreg/_03796_ ), .Z(\mreg/_00590_ ) );
MUX2_X1 \mreg/_10260_ ( .A(\mreg/_04142_ ), .B(\mreg/_04947_ ), .S(\mreg/_03796_ ), .Z(\mreg/_00591_ ) );
MUX2_X1 \mreg/_10261_ ( .A(\mreg/_04143_ ), .B(\mreg/_04948_ ), .S(\mreg/_03796_ ), .Z(\mreg/_00592_ ) );
MUX2_X1 \mreg/_10262_ ( .A(\mreg/_04144_ ), .B(\mreg/_04949_ ), .S(\mreg/_03796_ ), .Z(\mreg/_00593_ ) );
BUF_X4 \mreg/_10263_ ( .A(\mreg/_03794_ ), .Z(\mreg/_03797_ ) );
MUX2_X1 \mreg/_10264_ ( .A(\mreg/_04146_ ), .B(\mreg/_04951_ ), .S(\mreg/_03797_ ), .Z(\mreg/_00594_ ) );
MUX2_X1 \mreg/_10265_ ( .A(\mreg/_04147_ ), .B(\mreg/_04952_ ), .S(\mreg/_03797_ ), .Z(\mreg/_00595_ ) );
MUX2_X1 \mreg/_10266_ ( .A(\mreg/_04148_ ), .B(\mreg/_04953_ ), .S(\mreg/_03797_ ), .Z(\mreg/_00596_ ) );
MUX2_X1 \mreg/_10267_ ( .A(\mreg/_04149_ ), .B(\mreg/_04954_ ), .S(\mreg/_03797_ ), .Z(\mreg/_00597_ ) );
MUX2_X1 \mreg/_10268_ ( .A(\mreg/_04150_ ), .B(\mreg/_04955_ ), .S(\mreg/_03797_ ), .Z(\mreg/_00598_ ) );
MUX2_X1 \mreg/_10269_ ( .A(\mreg/_04151_ ), .B(\mreg/_04956_ ), .S(\mreg/_03797_ ), .Z(\mreg/_00599_ ) );
MUX2_X1 \mreg/_10270_ ( .A(\mreg/_04152_ ), .B(\mreg/_04957_ ), .S(\mreg/_03797_ ), .Z(\mreg/_00600_ ) );
MUX2_X1 \mreg/_10271_ ( .A(\mreg/_04153_ ), .B(\mreg/_04958_ ), .S(\mreg/_03797_ ), .Z(\mreg/_00601_ ) );
MUX2_X1 \mreg/_10272_ ( .A(\mreg/_04154_ ), .B(\mreg/_04959_ ), .S(\mreg/_03797_ ), .Z(\mreg/_00602_ ) );
MUX2_X1 \mreg/_10273_ ( .A(\mreg/_04155_ ), .B(\mreg/_04960_ ), .S(\mreg/_03797_ ), .Z(\mreg/_00603_ ) );
MUX2_X1 \mreg/_10274_ ( .A(\mreg/_04157_ ), .B(\mreg/_04962_ ), .S(\mreg/_03794_ ), .Z(\mreg/_00604_ ) );
MUX2_X1 \mreg/_10275_ ( .A(\mreg/_04158_ ), .B(\mreg/_04963_ ), .S(\mreg/_03794_ ), .Z(\mreg/_00605_ ) );
OR3_X1 \mreg/_10276_ ( .A1(\mreg/_03706_ ), .A2(\mreg/_03707_ ), .A3(\mreg/_03692_ ), .ZN(\mreg/_03798_ ) );
NOR2_X4 \mreg/_10277_ ( .A1(\mreg/_03798_ ), .A2(\mreg/_03783_ ), .ZN(\mreg/_03799_ ) );
BUF_X4 \mreg/_10278_ ( .A(\mreg/_03799_ ), .Z(\mreg/_03800_ ) );
MUX2_X1 \mreg/_10279_ ( .A(\mreg/_04166_ ), .B(\mreg/_04939_ ), .S(\mreg/_03800_ ), .Z(\mreg/_00606_ ) );
MUX2_X1 \mreg/_10280_ ( .A(\mreg/_04177_ ), .B(\mreg/_04950_ ), .S(\mreg/_03800_ ), .Z(\mreg/_00607_ ) );
MUX2_X1 \mreg/_10281_ ( .A(\mreg/_04188_ ), .B(\mreg/_04961_ ), .S(\mreg/_03800_ ), .Z(\mreg/_00608_ ) );
MUX2_X1 \mreg/_10282_ ( .A(\mreg/_04191_ ), .B(\mreg/_04964_ ), .S(\mreg/_03800_ ), .Z(\mreg/_00609_ ) );
MUX2_X1 \mreg/_10283_ ( .A(\mreg/_04192_ ), .B(\mreg/_04965_ ), .S(\mreg/_03800_ ), .Z(\mreg/_00610_ ) );
MUX2_X1 \mreg/_10284_ ( .A(\mreg/_04193_ ), .B(\mreg/_04966_ ), .S(\mreg/_03800_ ), .Z(\mreg/_00611_ ) );
MUX2_X1 \mreg/_10285_ ( .A(\mreg/_04194_ ), .B(\mreg/_04967_ ), .S(\mreg/_03800_ ), .Z(\mreg/_00612_ ) );
MUX2_X1 \mreg/_10286_ ( .A(\mreg/_04195_ ), .B(\mreg/_04968_ ), .S(\mreg/_03800_ ), .Z(\mreg/_00613_ ) );
MUX2_X1 \mreg/_10287_ ( .A(\mreg/_04196_ ), .B(\mreg/_04969_ ), .S(\mreg/_03800_ ), .Z(\mreg/_00614_ ) );
MUX2_X1 \mreg/_10288_ ( .A(\mreg/_04197_ ), .B(\mreg/_04970_ ), .S(\mreg/_03800_ ), .Z(\mreg/_00615_ ) );
BUF_X4 \mreg/_10289_ ( .A(\mreg/_03799_ ), .Z(\mreg/_03801_ ) );
MUX2_X1 \mreg/_10290_ ( .A(\mreg/_04167_ ), .B(\mreg/_04940_ ), .S(\mreg/_03801_ ), .Z(\mreg/_00616_ ) );
MUX2_X1 \mreg/_10291_ ( .A(\mreg/_04168_ ), .B(\mreg/_04941_ ), .S(\mreg/_03801_ ), .Z(\mreg/_00617_ ) );
MUX2_X1 \mreg/_10292_ ( .A(\mreg/_04169_ ), .B(\mreg/_04942_ ), .S(\mreg/_03801_ ), .Z(\mreg/_00618_ ) );
MUX2_X1 \mreg/_10293_ ( .A(\mreg/_04170_ ), .B(\mreg/_04943_ ), .S(\mreg/_03801_ ), .Z(\mreg/_00619_ ) );
MUX2_X1 \mreg/_10294_ ( .A(\mreg/_04171_ ), .B(\mreg/_04944_ ), .S(\mreg/_03801_ ), .Z(\mreg/_00620_ ) );
MUX2_X1 \mreg/_10295_ ( .A(\mreg/_04172_ ), .B(\mreg/_04945_ ), .S(\mreg/_03801_ ), .Z(\mreg/_00621_ ) );
MUX2_X1 \mreg/_10296_ ( .A(\mreg/_04173_ ), .B(\mreg/_04946_ ), .S(\mreg/_03801_ ), .Z(\mreg/_00622_ ) );
MUX2_X1 \mreg/_10297_ ( .A(\mreg/_04174_ ), .B(\mreg/_04947_ ), .S(\mreg/_03801_ ), .Z(\mreg/_00623_ ) );
MUX2_X1 \mreg/_10298_ ( .A(\mreg/_04175_ ), .B(\mreg/_04948_ ), .S(\mreg/_03801_ ), .Z(\mreg/_00624_ ) );
MUX2_X1 \mreg/_10299_ ( .A(\mreg/_04176_ ), .B(\mreg/_04949_ ), .S(\mreg/_03801_ ), .Z(\mreg/_00625_ ) );
BUF_X4 \mreg/_10300_ ( .A(\mreg/_03799_ ), .Z(\mreg/_03802_ ) );
MUX2_X1 \mreg/_10301_ ( .A(\mreg/_04178_ ), .B(\mreg/_04951_ ), .S(\mreg/_03802_ ), .Z(\mreg/_00626_ ) );
MUX2_X1 \mreg/_10302_ ( .A(\mreg/_04179_ ), .B(\mreg/_04952_ ), .S(\mreg/_03802_ ), .Z(\mreg/_00627_ ) );
MUX2_X1 \mreg/_10303_ ( .A(\mreg/_04180_ ), .B(\mreg/_04953_ ), .S(\mreg/_03802_ ), .Z(\mreg/_00628_ ) );
MUX2_X1 \mreg/_10304_ ( .A(\mreg/_04181_ ), .B(\mreg/_04954_ ), .S(\mreg/_03802_ ), .Z(\mreg/_00629_ ) );
MUX2_X1 \mreg/_10305_ ( .A(\mreg/_04182_ ), .B(\mreg/_04955_ ), .S(\mreg/_03802_ ), .Z(\mreg/_00630_ ) );
MUX2_X1 \mreg/_10306_ ( .A(\mreg/_04183_ ), .B(\mreg/_04956_ ), .S(\mreg/_03802_ ), .Z(\mreg/_00631_ ) );
MUX2_X1 \mreg/_10307_ ( .A(\mreg/_04184_ ), .B(\mreg/_04957_ ), .S(\mreg/_03802_ ), .Z(\mreg/_00632_ ) );
MUX2_X1 \mreg/_10308_ ( .A(\mreg/_04185_ ), .B(\mreg/_04958_ ), .S(\mreg/_03802_ ), .Z(\mreg/_00633_ ) );
MUX2_X1 \mreg/_10309_ ( .A(\mreg/_04186_ ), .B(\mreg/_04959_ ), .S(\mreg/_03802_ ), .Z(\mreg/_00634_ ) );
MUX2_X1 \mreg/_10310_ ( .A(\mreg/_04187_ ), .B(\mreg/_04960_ ), .S(\mreg/_03802_ ), .Z(\mreg/_00635_ ) );
MUX2_X1 \mreg/_10311_ ( .A(\mreg/_04189_ ), .B(\mreg/_04962_ ), .S(\mreg/_03799_ ), .Z(\mreg/_00636_ ) );
MUX2_X1 \mreg/_10312_ ( .A(\mreg/_04190_ ), .B(\mreg/_04963_ ), .S(\mreg/_03799_ ), .Z(\mreg/_00637_ ) );
NAND4_X1 \mreg/_10313_ ( .A1(\mreg/_03690_ ), .A2(\mreg/_04938_ ), .A3(\mreg/_03705_ ), .A4(\mreg/_04935_ ), .ZN(\mreg/_03803_ ) );
NOR2_X1 \mreg/_10314_ ( .A1(\mreg/_03696_ ), .A2(\mreg/_03803_ ), .ZN(\mreg/_03804_ ) );
BUF_X4 \mreg/_10315_ ( .A(\mreg/_03804_ ), .Z(\mreg/_03805_ ) );
MUX2_X1 \mreg/_10316_ ( .A(\mreg/_04198_ ), .B(\mreg/_04939_ ), .S(\mreg/_03805_ ), .Z(\mreg/_00638_ ) );
MUX2_X1 \mreg/_10317_ ( .A(\mreg/_04209_ ), .B(\mreg/_04950_ ), .S(\mreg/_03805_ ), .Z(\mreg/_00639_ ) );
MUX2_X1 \mreg/_10318_ ( .A(\mreg/_04220_ ), .B(\mreg/_04961_ ), .S(\mreg/_03805_ ), .Z(\mreg/_00640_ ) );
MUX2_X1 \mreg/_10319_ ( .A(\mreg/_04223_ ), .B(\mreg/_04964_ ), .S(\mreg/_03805_ ), .Z(\mreg/_00641_ ) );
MUX2_X1 \mreg/_10320_ ( .A(\mreg/_04224_ ), .B(\mreg/_04965_ ), .S(\mreg/_03805_ ), .Z(\mreg/_00642_ ) );
MUX2_X1 \mreg/_10321_ ( .A(\mreg/_04225_ ), .B(\mreg/_04966_ ), .S(\mreg/_03805_ ), .Z(\mreg/_00643_ ) );
MUX2_X1 \mreg/_10322_ ( .A(\mreg/_04226_ ), .B(\mreg/_04967_ ), .S(\mreg/_03805_ ), .Z(\mreg/_00644_ ) );
MUX2_X1 \mreg/_10323_ ( .A(\mreg/_04227_ ), .B(\mreg/_04968_ ), .S(\mreg/_03805_ ), .Z(\mreg/_00645_ ) );
MUX2_X1 \mreg/_10324_ ( .A(\mreg/_04228_ ), .B(\mreg/_04969_ ), .S(\mreg/_03805_ ), .Z(\mreg/_00646_ ) );
MUX2_X1 \mreg/_10325_ ( .A(\mreg/_04229_ ), .B(\mreg/_04970_ ), .S(\mreg/_03805_ ), .Z(\mreg/_00647_ ) );
BUF_X4 \mreg/_10326_ ( .A(\mreg/_03804_ ), .Z(\mreg/_03806_ ) );
MUX2_X1 \mreg/_10327_ ( .A(\mreg/_04199_ ), .B(\mreg/_04940_ ), .S(\mreg/_03806_ ), .Z(\mreg/_00648_ ) );
MUX2_X1 \mreg/_10328_ ( .A(\mreg/_04200_ ), .B(\mreg/_04941_ ), .S(\mreg/_03806_ ), .Z(\mreg/_00649_ ) );
MUX2_X1 \mreg/_10329_ ( .A(\mreg/_04201_ ), .B(\mreg/_04942_ ), .S(\mreg/_03806_ ), .Z(\mreg/_00650_ ) );
MUX2_X1 \mreg/_10330_ ( .A(\mreg/_04202_ ), .B(\mreg/_04943_ ), .S(\mreg/_03806_ ), .Z(\mreg/_00651_ ) );
MUX2_X1 \mreg/_10331_ ( .A(\mreg/_04203_ ), .B(\mreg/_04944_ ), .S(\mreg/_03806_ ), .Z(\mreg/_00652_ ) );
MUX2_X1 \mreg/_10332_ ( .A(\mreg/_04204_ ), .B(\mreg/_04945_ ), .S(\mreg/_03806_ ), .Z(\mreg/_00653_ ) );
MUX2_X1 \mreg/_10333_ ( .A(\mreg/_04205_ ), .B(\mreg/_04946_ ), .S(\mreg/_03806_ ), .Z(\mreg/_00654_ ) );
MUX2_X1 \mreg/_10334_ ( .A(\mreg/_04206_ ), .B(\mreg/_04947_ ), .S(\mreg/_03806_ ), .Z(\mreg/_00655_ ) );
MUX2_X1 \mreg/_10335_ ( .A(\mreg/_04207_ ), .B(\mreg/_04948_ ), .S(\mreg/_03806_ ), .Z(\mreg/_00656_ ) );
MUX2_X1 \mreg/_10336_ ( .A(\mreg/_04208_ ), .B(\mreg/_04949_ ), .S(\mreg/_03806_ ), .Z(\mreg/_00657_ ) );
BUF_X4 \mreg/_10337_ ( .A(\mreg/_03804_ ), .Z(\mreg/_03807_ ) );
MUX2_X1 \mreg/_10338_ ( .A(\mreg/_04210_ ), .B(\mreg/_04951_ ), .S(\mreg/_03807_ ), .Z(\mreg/_00658_ ) );
MUX2_X1 \mreg/_10339_ ( .A(\mreg/_04211_ ), .B(\mreg/_04952_ ), .S(\mreg/_03807_ ), .Z(\mreg/_00659_ ) );
MUX2_X1 \mreg/_10340_ ( .A(\mreg/_04212_ ), .B(\mreg/_04953_ ), .S(\mreg/_03807_ ), .Z(\mreg/_00660_ ) );
MUX2_X1 \mreg/_10341_ ( .A(\mreg/_04213_ ), .B(\mreg/_04954_ ), .S(\mreg/_03807_ ), .Z(\mreg/_00661_ ) );
MUX2_X1 \mreg/_10342_ ( .A(\mreg/_04214_ ), .B(\mreg/_04955_ ), .S(\mreg/_03807_ ), .Z(\mreg/_00662_ ) );
MUX2_X1 \mreg/_10343_ ( .A(\mreg/_04215_ ), .B(\mreg/_04956_ ), .S(\mreg/_03807_ ), .Z(\mreg/_00663_ ) );
MUX2_X1 \mreg/_10344_ ( .A(\mreg/_04216_ ), .B(\mreg/_04957_ ), .S(\mreg/_03807_ ), .Z(\mreg/_00664_ ) );
MUX2_X1 \mreg/_10345_ ( .A(\mreg/_04217_ ), .B(\mreg/_04958_ ), .S(\mreg/_03807_ ), .Z(\mreg/_00665_ ) );
MUX2_X1 \mreg/_10346_ ( .A(\mreg/_04218_ ), .B(\mreg/_04959_ ), .S(\mreg/_03807_ ), .Z(\mreg/_00666_ ) );
MUX2_X1 \mreg/_10347_ ( .A(\mreg/_04219_ ), .B(\mreg/_04960_ ), .S(\mreg/_03807_ ), .Z(\mreg/_00667_ ) );
MUX2_X1 \mreg/_10348_ ( .A(\mreg/_04221_ ), .B(\mreg/_04962_ ), .S(\mreg/_03804_ ), .Z(\mreg/_00668_ ) );
MUX2_X1 \mreg/_10349_ ( .A(\mreg/_04222_ ), .B(\mreg/_04963_ ), .S(\mreg/_03804_ ), .Z(\mreg/_00669_ ) );
NAND4_X1 \mreg/_10350_ ( .A1(\mreg/_03690_ ), .A2(\mreg/_04938_ ), .A3(\mreg/_04934_ ), .A4(\mreg/_04935_ ), .ZN(\mreg/_03808_ ) );
NOR2_X1 \mreg/_10351_ ( .A1(\mreg/_03696_ ), .A2(\mreg/_03808_ ), .ZN(\mreg/_03809_ ) );
BUF_X4 \mreg/_10352_ ( .A(\mreg/_03809_ ), .Z(\mreg/_03810_ ) );
MUX2_X1 \mreg/_10353_ ( .A(\mreg/_04230_ ), .B(\mreg/_04939_ ), .S(\mreg/_03810_ ), .Z(\mreg/_00670_ ) );
MUX2_X1 \mreg/_10354_ ( .A(\mreg/_04241_ ), .B(\mreg/_04950_ ), .S(\mreg/_03810_ ), .Z(\mreg/_00671_ ) );
MUX2_X1 \mreg/_10355_ ( .A(\mreg/_04252_ ), .B(\mreg/_04961_ ), .S(\mreg/_03810_ ), .Z(\mreg/_00672_ ) );
MUX2_X1 \mreg/_10356_ ( .A(\mreg/_04255_ ), .B(\mreg/_04964_ ), .S(\mreg/_03810_ ), .Z(\mreg/_00673_ ) );
MUX2_X1 \mreg/_10357_ ( .A(\mreg/_04256_ ), .B(\mreg/_04965_ ), .S(\mreg/_03810_ ), .Z(\mreg/_00674_ ) );
MUX2_X1 \mreg/_10358_ ( .A(\mreg/_04257_ ), .B(\mreg/_04966_ ), .S(\mreg/_03810_ ), .Z(\mreg/_00675_ ) );
MUX2_X1 \mreg/_10359_ ( .A(\mreg/_04258_ ), .B(\mreg/_04967_ ), .S(\mreg/_03810_ ), .Z(\mreg/_00676_ ) );
MUX2_X1 \mreg/_10360_ ( .A(\mreg/_04259_ ), .B(\mreg/_04968_ ), .S(\mreg/_03810_ ), .Z(\mreg/_00677_ ) );
MUX2_X1 \mreg/_10361_ ( .A(\mreg/_04260_ ), .B(\mreg/_04969_ ), .S(\mreg/_03810_ ), .Z(\mreg/_00678_ ) );
MUX2_X1 \mreg/_10362_ ( .A(\mreg/_04261_ ), .B(\mreg/_04970_ ), .S(\mreg/_03810_ ), .Z(\mreg/_00679_ ) );
BUF_X4 \mreg/_10363_ ( .A(\mreg/_03809_ ), .Z(\mreg/_03811_ ) );
MUX2_X1 \mreg/_10364_ ( .A(\mreg/_04231_ ), .B(\mreg/_04940_ ), .S(\mreg/_03811_ ), .Z(\mreg/_00680_ ) );
MUX2_X1 \mreg/_10365_ ( .A(\mreg/_04232_ ), .B(\mreg/_04941_ ), .S(\mreg/_03811_ ), .Z(\mreg/_00681_ ) );
MUX2_X1 \mreg/_10366_ ( .A(\mreg/_04233_ ), .B(\mreg/_04942_ ), .S(\mreg/_03811_ ), .Z(\mreg/_00682_ ) );
MUX2_X1 \mreg/_10367_ ( .A(\mreg/_04234_ ), .B(\mreg/_04943_ ), .S(\mreg/_03811_ ), .Z(\mreg/_00683_ ) );
MUX2_X1 \mreg/_10368_ ( .A(\mreg/_04235_ ), .B(\mreg/_04944_ ), .S(\mreg/_03811_ ), .Z(\mreg/_00684_ ) );
MUX2_X1 \mreg/_10369_ ( .A(\mreg/_04236_ ), .B(\mreg/_04945_ ), .S(\mreg/_03811_ ), .Z(\mreg/_00685_ ) );
MUX2_X1 \mreg/_10370_ ( .A(\mreg/_04237_ ), .B(\mreg/_04946_ ), .S(\mreg/_03811_ ), .Z(\mreg/_00686_ ) );
MUX2_X1 \mreg/_10371_ ( .A(\mreg/_04238_ ), .B(\mreg/_04947_ ), .S(\mreg/_03811_ ), .Z(\mreg/_00687_ ) );
MUX2_X1 \mreg/_10372_ ( .A(\mreg/_04239_ ), .B(\mreg/_04948_ ), .S(\mreg/_03811_ ), .Z(\mreg/_00688_ ) );
MUX2_X1 \mreg/_10373_ ( .A(\mreg/_04240_ ), .B(\mreg/_04949_ ), .S(\mreg/_03811_ ), .Z(\mreg/_00689_ ) );
BUF_X4 \mreg/_10374_ ( .A(\mreg/_03809_ ), .Z(\mreg/_03812_ ) );
MUX2_X1 \mreg/_10375_ ( .A(\mreg/_04242_ ), .B(\mreg/_04951_ ), .S(\mreg/_03812_ ), .Z(\mreg/_00690_ ) );
MUX2_X1 \mreg/_10376_ ( .A(\mreg/_04243_ ), .B(\mreg/_04952_ ), .S(\mreg/_03812_ ), .Z(\mreg/_00691_ ) );
MUX2_X1 \mreg/_10377_ ( .A(\mreg/_04244_ ), .B(\mreg/_04953_ ), .S(\mreg/_03812_ ), .Z(\mreg/_00692_ ) );
MUX2_X1 \mreg/_10378_ ( .A(\mreg/_04245_ ), .B(\mreg/_04954_ ), .S(\mreg/_03812_ ), .Z(\mreg/_00693_ ) );
MUX2_X1 \mreg/_10379_ ( .A(\mreg/_04246_ ), .B(\mreg/_04955_ ), .S(\mreg/_03812_ ), .Z(\mreg/_00694_ ) );
MUX2_X1 \mreg/_10380_ ( .A(\mreg/_04247_ ), .B(\mreg/_04956_ ), .S(\mreg/_03812_ ), .Z(\mreg/_00695_ ) );
MUX2_X1 \mreg/_10381_ ( .A(\mreg/_04248_ ), .B(\mreg/_04957_ ), .S(\mreg/_03812_ ), .Z(\mreg/_00696_ ) );
MUX2_X1 \mreg/_10382_ ( .A(\mreg/_04249_ ), .B(\mreg/_04958_ ), .S(\mreg/_03812_ ), .Z(\mreg/_00697_ ) );
MUX2_X1 \mreg/_10383_ ( .A(\mreg/_04250_ ), .B(\mreg/_04959_ ), .S(\mreg/_03812_ ), .Z(\mreg/_00698_ ) );
MUX2_X1 \mreg/_10384_ ( .A(\mreg/_04251_ ), .B(\mreg/_04960_ ), .S(\mreg/_03812_ ), .Z(\mreg/_00699_ ) );
MUX2_X1 \mreg/_10385_ ( .A(\mreg/_04253_ ), .B(\mreg/_04962_ ), .S(\mreg/_03809_ ), .Z(\mreg/_00700_ ) );
MUX2_X1 \mreg/_10386_ ( .A(\mreg/_04254_ ), .B(\mreg/_04963_ ), .S(\mreg/_03809_ ), .Z(\mreg/_00701_ ) );
OR3_X1 \mreg/_10387_ ( .A1(\mreg/_03726_ ), .A2(\mreg/_03727_ ), .A3(\mreg/_03692_ ), .ZN(\mreg/_03813_ ) );
NOR2_X4 \mreg/_10388_ ( .A1(\mreg/_03813_ ), .A2(\mreg/_03783_ ), .ZN(\mreg/_03814_ ) );
BUF_X4 \mreg/_10389_ ( .A(\mreg/_03814_ ), .Z(\mreg/_03815_ ) );
MUX2_X1 \mreg/_10390_ ( .A(\mreg/_04294_ ), .B(\mreg/_04939_ ), .S(\mreg/_03815_ ), .Z(\mreg/_00702_ ) );
MUX2_X1 \mreg/_10391_ ( .A(\mreg/_04305_ ), .B(\mreg/_04950_ ), .S(\mreg/_03815_ ), .Z(\mreg/_00703_ ) );
MUX2_X1 \mreg/_10392_ ( .A(\mreg/_04316_ ), .B(\mreg/_04961_ ), .S(\mreg/_03815_ ), .Z(\mreg/_00704_ ) );
MUX2_X1 \mreg/_10393_ ( .A(\mreg/_04319_ ), .B(\mreg/_04964_ ), .S(\mreg/_03815_ ), .Z(\mreg/_00705_ ) );
MUX2_X1 \mreg/_10394_ ( .A(\mreg/_04320_ ), .B(\mreg/_04965_ ), .S(\mreg/_03815_ ), .Z(\mreg/_00706_ ) );
MUX2_X1 \mreg/_10395_ ( .A(\mreg/_04321_ ), .B(\mreg/_04966_ ), .S(\mreg/_03815_ ), .Z(\mreg/_00707_ ) );
MUX2_X1 \mreg/_10396_ ( .A(\mreg/_04322_ ), .B(\mreg/_04967_ ), .S(\mreg/_03815_ ), .Z(\mreg/_00708_ ) );
MUX2_X1 \mreg/_10397_ ( .A(\mreg/_04323_ ), .B(\mreg/_04968_ ), .S(\mreg/_03815_ ), .Z(\mreg/_00709_ ) );
MUX2_X1 \mreg/_10398_ ( .A(\mreg/_04324_ ), .B(\mreg/_04969_ ), .S(\mreg/_03815_ ), .Z(\mreg/_00710_ ) );
MUX2_X1 \mreg/_10399_ ( .A(\mreg/_04325_ ), .B(\mreg/_04970_ ), .S(\mreg/_03815_ ), .Z(\mreg/_00711_ ) );
BUF_X4 \mreg/_10400_ ( .A(\mreg/_03814_ ), .Z(\mreg/_03816_ ) );
MUX2_X1 \mreg/_10401_ ( .A(\mreg/_04295_ ), .B(\mreg/_04940_ ), .S(\mreg/_03816_ ), .Z(\mreg/_00712_ ) );
MUX2_X1 \mreg/_10402_ ( .A(\mreg/_04296_ ), .B(\mreg/_04941_ ), .S(\mreg/_03816_ ), .Z(\mreg/_00713_ ) );
MUX2_X1 \mreg/_10403_ ( .A(\mreg/_04297_ ), .B(\mreg/_04942_ ), .S(\mreg/_03816_ ), .Z(\mreg/_00714_ ) );
MUX2_X1 \mreg/_10404_ ( .A(\mreg/_04298_ ), .B(\mreg/_04943_ ), .S(\mreg/_03816_ ), .Z(\mreg/_00715_ ) );
MUX2_X1 \mreg/_10405_ ( .A(\mreg/_04299_ ), .B(\mreg/_04944_ ), .S(\mreg/_03816_ ), .Z(\mreg/_00716_ ) );
MUX2_X1 \mreg/_10406_ ( .A(\mreg/_04300_ ), .B(\mreg/_04945_ ), .S(\mreg/_03816_ ), .Z(\mreg/_00717_ ) );
MUX2_X1 \mreg/_10407_ ( .A(\mreg/_04301_ ), .B(\mreg/_04946_ ), .S(\mreg/_03816_ ), .Z(\mreg/_00718_ ) );
MUX2_X1 \mreg/_10408_ ( .A(\mreg/_04302_ ), .B(\mreg/_04947_ ), .S(\mreg/_03816_ ), .Z(\mreg/_00719_ ) );
MUX2_X1 \mreg/_10409_ ( .A(\mreg/_04303_ ), .B(\mreg/_04948_ ), .S(\mreg/_03816_ ), .Z(\mreg/_00720_ ) );
MUX2_X1 \mreg/_10410_ ( .A(\mreg/_04304_ ), .B(\mreg/_04949_ ), .S(\mreg/_03816_ ), .Z(\mreg/_00721_ ) );
BUF_X4 \mreg/_10411_ ( .A(\mreg/_03814_ ), .Z(\mreg/_03817_ ) );
MUX2_X1 \mreg/_10412_ ( .A(\mreg/_04306_ ), .B(\mreg/_04951_ ), .S(\mreg/_03817_ ), .Z(\mreg/_00722_ ) );
MUX2_X1 \mreg/_10413_ ( .A(\mreg/_04307_ ), .B(\mreg/_04952_ ), .S(\mreg/_03817_ ), .Z(\mreg/_00723_ ) );
MUX2_X1 \mreg/_10414_ ( .A(\mreg/_04308_ ), .B(\mreg/_04953_ ), .S(\mreg/_03817_ ), .Z(\mreg/_00724_ ) );
MUX2_X1 \mreg/_10415_ ( .A(\mreg/_04309_ ), .B(\mreg/_04954_ ), .S(\mreg/_03817_ ), .Z(\mreg/_00725_ ) );
MUX2_X1 \mreg/_10416_ ( .A(\mreg/_04310_ ), .B(\mreg/_04955_ ), .S(\mreg/_03817_ ), .Z(\mreg/_00726_ ) );
MUX2_X1 \mreg/_10417_ ( .A(\mreg/_04311_ ), .B(\mreg/_04956_ ), .S(\mreg/_03817_ ), .Z(\mreg/_00727_ ) );
MUX2_X1 \mreg/_10418_ ( .A(\mreg/_04312_ ), .B(\mreg/_04957_ ), .S(\mreg/_03817_ ), .Z(\mreg/_00728_ ) );
MUX2_X1 \mreg/_10419_ ( .A(\mreg/_04313_ ), .B(\mreg/_04958_ ), .S(\mreg/_03817_ ), .Z(\mreg/_00729_ ) );
MUX2_X1 \mreg/_10420_ ( .A(\mreg/_04314_ ), .B(\mreg/_04959_ ), .S(\mreg/_03817_ ), .Z(\mreg/_00730_ ) );
MUX2_X1 \mreg/_10421_ ( .A(\mreg/_04315_ ), .B(\mreg/_04960_ ), .S(\mreg/_03817_ ), .Z(\mreg/_00731_ ) );
MUX2_X1 \mreg/_10422_ ( .A(\mreg/_04317_ ), .B(\mreg/_04962_ ), .S(\mreg/_03814_ ), .Z(\mreg/_00732_ ) );
MUX2_X1 \mreg/_10423_ ( .A(\mreg/_04318_ ), .B(\mreg/_04963_ ), .S(\mreg/_03814_ ), .Z(\mreg/_00733_ ) );
NAND2_X1 \mreg/_10424_ ( .A1(\mreg/_03733_ ), .A2(\mreg/_04938_ ), .ZN(\mreg/_03818_ ) );
NOR2_X1 \mreg/_10425_ ( .A1(\mreg/_03818_ ), .A2(\mreg/_03783_ ), .ZN(\mreg/_03819_ ) );
BUF_X4 \mreg/_10426_ ( .A(\mreg/_03819_ ), .Z(\mreg/_03820_ ) );
MUX2_X1 \mreg/_10427_ ( .A(\mreg/_04326_ ), .B(\mreg/_04939_ ), .S(\mreg/_03820_ ), .Z(\mreg/_00734_ ) );
MUX2_X1 \mreg/_10428_ ( .A(\mreg/_04337_ ), .B(\mreg/_04950_ ), .S(\mreg/_03820_ ), .Z(\mreg/_00735_ ) );
MUX2_X1 \mreg/_10429_ ( .A(\mreg/_04348_ ), .B(\mreg/_04961_ ), .S(\mreg/_03820_ ), .Z(\mreg/_00736_ ) );
MUX2_X1 \mreg/_10430_ ( .A(\mreg/_04351_ ), .B(\mreg/_04964_ ), .S(\mreg/_03820_ ), .Z(\mreg/_00737_ ) );
MUX2_X1 \mreg/_10431_ ( .A(\mreg/_04352_ ), .B(\mreg/_04965_ ), .S(\mreg/_03820_ ), .Z(\mreg/_00738_ ) );
MUX2_X1 \mreg/_10432_ ( .A(\mreg/_04353_ ), .B(\mreg/_04966_ ), .S(\mreg/_03820_ ), .Z(\mreg/_00739_ ) );
MUX2_X1 \mreg/_10433_ ( .A(\mreg/_04354_ ), .B(\mreg/_04967_ ), .S(\mreg/_03820_ ), .Z(\mreg/_00740_ ) );
MUX2_X1 \mreg/_10434_ ( .A(\mreg/_04355_ ), .B(\mreg/_04968_ ), .S(\mreg/_03820_ ), .Z(\mreg/_00741_ ) );
MUX2_X1 \mreg/_10435_ ( .A(\mreg/_04356_ ), .B(\mreg/_04969_ ), .S(\mreg/_03820_ ), .Z(\mreg/_00742_ ) );
MUX2_X1 \mreg/_10436_ ( .A(\mreg/_04357_ ), .B(\mreg/_04970_ ), .S(\mreg/_03820_ ), .Z(\mreg/_00743_ ) );
BUF_X4 \mreg/_10437_ ( .A(\mreg/_03819_ ), .Z(\mreg/_03821_ ) );
MUX2_X1 \mreg/_10438_ ( .A(\mreg/_04327_ ), .B(\mreg/_04940_ ), .S(\mreg/_03821_ ), .Z(\mreg/_00744_ ) );
MUX2_X1 \mreg/_10439_ ( .A(\mreg/_04328_ ), .B(\mreg/_04941_ ), .S(\mreg/_03821_ ), .Z(\mreg/_00745_ ) );
MUX2_X1 \mreg/_10440_ ( .A(\mreg/_04329_ ), .B(\mreg/_04942_ ), .S(\mreg/_03821_ ), .Z(\mreg/_00746_ ) );
MUX2_X1 \mreg/_10441_ ( .A(\mreg/_04330_ ), .B(\mreg/_04943_ ), .S(\mreg/_03821_ ), .Z(\mreg/_00747_ ) );
MUX2_X1 \mreg/_10442_ ( .A(\mreg/_04331_ ), .B(\mreg/_04944_ ), .S(\mreg/_03821_ ), .Z(\mreg/_00748_ ) );
MUX2_X1 \mreg/_10443_ ( .A(\mreg/_04332_ ), .B(\mreg/_04945_ ), .S(\mreg/_03821_ ), .Z(\mreg/_00749_ ) );
MUX2_X1 \mreg/_10444_ ( .A(\mreg/_04333_ ), .B(\mreg/_04946_ ), .S(\mreg/_03821_ ), .Z(\mreg/_00750_ ) );
MUX2_X1 \mreg/_10445_ ( .A(\mreg/_04334_ ), .B(\mreg/_04947_ ), .S(\mreg/_03821_ ), .Z(\mreg/_00751_ ) );
MUX2_X1 \mreg/_10446_ ( .A(\mreg/_04335_ ), .B(\mreg/_04948_ ), .S(\mreg/_03821_ ), .Z(\mreg/_00752_ ) );
MUX2_X1 \mreg/_10447_ ( .A(\mreg/_04336_ ), .B(\mreg/_04949_ ), .S(\mreg/_03821_ ), .Z(\mreg/_00753_ ) );
BUF_X4 \mreg/_10448_ ( .A(\mreg/_03819_ ), .Z(\mreg/_03822_ ) );
MUX2_X1 \mreg/_10449_ ( .A(\mreg/_04338_ ), .B(\mreg/_04951_ ), .S(\mreg/_03822_ ), .Z(\mreg/_00754_ ) );
MUX2_X1 \mreg/_10450_ ( .A(\mreg/_04339_ ), .B(\mreg/_04952_ ), .S(\mreg/_03822_ ), .Z(\mreg/_00755_ ) );
MUX2_X1 \mreg/_10451_ ( .A(\mreg/_04340_ ), .B(\mreg/_04953_ ), .S(\mreg/_03822_ ), .Z(\mreg/_00756_ ) );
MUX2_X1 \mreg/_10452_ ( .A(\mreg/_04341_ ), .B(\mreg/_04954_ ), .S(\mreg/_03822_ ), .Z(\mreg/_00757_ ) );
MUX2_X1 \mreg/_10453_ ( .A(\mreg/_04342_ ), .B(\mreg/_04955_ ), .S(\mreg/_03822_ ), .Z(\mreg/_00758_ ) );
MUX2_X1 \mreg/_10454_ ( .A(\mreg/_04343_ ), .B(\mreg/_04956_ ), .S(\mreg/_03822_ ), .Z(\mreg/_00759_ ) );
MUX2_X1 \mreg/_10455_ ( .A(\mreg/_04344_ ), .B(\mreg/_04957_ ), .S(\mreg/_03822_ ), .Z(\mreg/_00760_ ) );
MUX2_X1 \mreg/_10456_ ( .A(\mreg/_04345_ ), .B(\mreg/_04958_ ), .S(\mreg/_03822_ ), .Z(\mreg/_00761_ ) );
MUX2_X1 \mreg/_10457_ ( .A(\mreg/_04346_ ), .B(\mreg/_04959_ ), .S(\mreg/_03822_ ), .Z(\mreg/_00762_ ) );
MUX2_X1 \mreg/_10458_ ( .A(\mreg/_04347_ ), .B(\mreg/_04960_ ), .S(\mreg/_03822_ ), .Z(\mreg/_00763_ ) );
MUX2_X1 \mreg/_10459_ ( .A(\mreg/_04349_ ), .B(\mreg/_04962_ ), .S(\mreg/_03819_ ), .Z(\mreg/_00764_ ) );
MUX2_X1 \mreg/_10460_ ( .A(\mreg/_04350_ ), .B(\mreg/_04963_ ), .S(\mreg/_03819_ ), .Z(\mreg/_00765_ ) );
OR3_X1 \mreg/_10461_ ( .A1(\mreg/_03726_ ), .A2(\mreg/_03714_ ), .A3(\mreg/_03739_ ), .ZN(\mreg/_03823_ ) );
NOR2_X1 \mreg/_10462_ ( .A1(\mreg/_03823_ ), .A2(\mreg/_03783_ ), .ZN(\mreg/_03824_ ) );
BUF_X4 \mreg/_10463_ ( .A(\mreg/_03824_ ), .Z(\mreg/_03825_ ) );
MUX2_X1 \mreg/_10464_ ( .A(\mreg/_04358_ ), .B(\mreg/_04939_ ), .S(\mreg/_03825_ ), .Z(\mreg/_00766_ ) );
MUX2_X1 \mreg/_10465_ ( .A(\mreg/_04369_ ), .B(\mreg/_04950_ ), .S(\mreg/_03825_ ), .Z(\mreg/_00767_ ) );
MUX2_X1 \mreg/_10466_ ( .A(\mreg/_04380_ ), .B(\mreg/_04961_ ), .S(\mreg/_03825_ ), .Z(\mreg/_00768_ ) );
MUX2_X1 \mreg/_10467_ ( .A(\mreg/_04383_ ), .B(\mreg/_04964_ ), .S(\mreg/_03825_ ), .Z(\mreg/_00769_ ) );
MUX2_X1 \mreg/_10468_ ( .A(\mreg/_04384_ ), .B(\mreg/_04965_ ), .S(\mreg/_03825_ ), .Z(\mreg/_00770_ ) );
MUX2_X1 \mreg/_10469_ ( .A(\mreg/_04385_ ), .B(\mreg/_04966_ ), .S(\mreg/_03825_ ), .Z(\mreg/_00771_ ) );
MUX2_X1 \mreg/_10470_ ( .A(\mreg/_04386_ ), .B(\mreg/_04967_ ), .S(\mreg/_03825_ ), .Z(\mreg/_00772_ ) );
MUX2_X1 \mreg/_10471_ ( .A(\mreg/_04387_ ), .B(\mreg/_04968_ ), .S(\mreg/_03825_ ), .Z(\mreg/_00773_ ) );
MUX2_X1 \mreg/_10472_ ( .A(\mreg/_04388_ ), .B(\mreg/_04969_ ), .S(\mreg/_03825_ ), .Z(\mreg/_00774_ ) );
MUX2_X1 \mreg/_10473_ ( .A(\mreg/_04389_ ), .B(\mreg/_04970_ ), .S(\mreg/_03825_ ), .Z(\mreg/_00775_ ) );
BUF_X4 \mreg/_10474_ ( .A(\mreg/_03824_ ), .Z(\mreg/_03826_ ) );
MUX2_X1 \mreg/_10475_ ( .A(\mreg/_04359_ ), .B(\mreg/_04940_ ), .S(\mreg/_03826_ ), .Z(\mreg/_00776_ ) );
MUX2_X1 \mreg/_10476_ ( .A(\mreg/_04360_ ), .B(\mreg/_04941_ ), .S(\mreg/_03826_ ), .Z(\mreg/_00777_ ) );
MUX2_X1 \mreg/_10477_ ( .A(\mreg/_04361_ ), .B(\mreg/_04942_ ), .S(\mreg/_03826_ ), .Z(\mreg/_00778_ ) );
MUX2_X1 \mreg/_10478_ ( .A(\mreg/_04362_ ), .B(\mreg/_04943_ ), .S(\mreg/_03826_ ), .Z(\mreg/_00779_ ) );
MUX2_X1 \mreg/_10479_ ( .A(\mreg/_04363_ ), .B(\mreg/_04944_ ), .S(\mreg/_03826_ ), .Z(\mreg/_00780_ ) );
MUX2_X1 \mreg/_10480_ ( .A(\mreg/_04364_ ), .B(\mreg/_04945_ ), .S(\mreg/_03826_ ), .Z(\mreg/_00781_ ) );
MUX2_X1 \mreg/_10481_ ( .A(\mreg/_04365_ ), .B(\mreg/_04946_ ), .S(\mreg/_03826_ ), .Z(\mreg/_00782_ ) );
MUX2_X1 \mreg/_10482_ ( .A(\mreg/_04366_ ), .B(\mreg/_04947_ ), .S(\mreg/_03826_ ), .Z(\mreg/_00783_ ) );
MUX2_X1 \mreg/_10483_ ( .A(\mreg/_04367_ ), .B(\mreg/_04948_ ), .S(\mreg/_03826_ ), .Z(\mreg/_00784_ ) );
MUX2_X1 \mreg/_10484_ ( .A(\mreg/_04368_ ), .B(\mreg/_04949_ ), .S(\mreg/_03826_ ), .Z(\mreg/_00785_ ) );
BUF_X4 \mreg/_10485_ ( .A(\mreg/_03824_ ), .Z(\mreg/_03827_ ) );
MUX2_X1 \mreg/_10486_ ( .A(\mreg/_04370_ ), .B(\mreg/_04951_ ), .S(\mreg/_03827_ ), .Z(\mreg/_00786_ ) );
MUX2_X1 \mreg/_10487_ ( .A(\mreg/_04371_ ), .B(\mreg/_04952_ ), .S(\mreg/_03827_ ), .Z(\mreg/_00787_ ) );
MUX2_X1 \mreg/_10488_ ( .A(\mreg/_04372_ ), .B(\mreg/_04953_ ), .S(\mreg/_03827_ ), .Z(\mreg/_00788_ ) );
MUX2_X1 \mreg/_10489_ ( .A(\mreg/_04373_ ), .B(\mreg/_04954_ ), .S(\mreg/_03827_ ), .Z(\mreg/_00789_ ) );
MUX2_X1 \mreg/_10490_ ( .A(\mreg/_04374_ ), .B(\mreg/_04955_ ), .S(\mreg/_03827_ ), .Z(\mreg/_00790_ ) );
MUX2_X1 \mreg/_10491_ ( .A(\mreg/_04375_ ), .B(\mreg/_04956_ ), .S(\mreg/_03827_ ), .Z(\mreg/_00791_ ) );
MUX2_X1 \mreg/_10492_ ( .A(\mreg/_04376_ ), .B(\mreg/_04957_ ), .S(\mreg/_03827_ ), .Z(\mreg/_00792_ ) );
MUX2_X1 \mreg/_10493_ ( .A(\mreg/_04377_ ), .B(\mreg/_04958_ ), .S(\mreg/_03827_ ), .Z(\mreg/_00793_ ) );
MUX2_X1 \mreg/_10494_ ( .A(\mreg/_04378_ ), .B(\mreg/_04959_ ), .S(\mreg/_03827_ ), .Z(\mreg/_00794_ ) );
MUX2_X1 \mreg/_10495_ ( .A(\mreg/_04379_ ), .B(\mreg/_04960_ ), .S(\mreg/_03827_ ), .Z(\mreg/_00795_ ) );
MUX2_X1 \mreg/_10496_ ( .A(\mreg/_04381_ ), .B(\mreg/_04962_ ), .S(\mreg/_03824_ ), .Z(\mreg/_00796_ ) );
MUX2_X1 \mreg/_10497_ ( .A(\mreg/_04382_ ), .B(\mreg/_04963_ ), .S(\mreg/_03824_ ), .Z(\mreg/_00797_ ) );
OR4_X1 \mreg/_10498_ ( .A1(\mreg/_03692_ ), .A2(\mreg/_03698_ ), .A3(\mreg/_03725_ ), .A4(\mreg/_04937_ ), .ZN(\mreg/_03828_ ) );
NOR2_X1 \mreg/_10499_ ( .A1(\mreg/_03828_ ), .A2(\mreg/_03783_ ), .ZN(\mreg/_03829_ ) );
BUF_X4 \mreg/_10500_ ( .A(\mreg/_03829_ ), .Z(\mreg/_03830_ ) );
MUX2_X1 \mreg/_10501_ ( .A(\mreg/_04390_ ), .B(\mreg/_04939_ ), .S(\mreg/_03830_ ), .Z(\mreg/_00798_ ) );
MUX2_X1 \mreg/_10502_ ( .A(\mreg/_04401_ ), .B(\mreg/_04950_ ), .S(\mreg/_03830_ ), .Z(\mreg/_00799_ ) );
MUX2_X1 \mreg/_10503_ ( .A(\mreg/_04412_ ), .B(\mreg/_04961_ ), .S(\mreg/_03830_ ), .Z(\mreg/_00800_ ) );
MUX2_X1 \mreg/_10504_ ( .A(\mreg/_04415_ ), .B(\mreg/_04964_ ), .S(\mreg/_03830_ ), .Z(\mreg/_00801_ ) );
MUX2_X1 \mreg/_10505_ ( .A(\mreg/_04416_ ), .B(\mreg/_04965_ ), .S(\mreg/_03830_ ), .Z(\mreg/_00802_ ) );
MUX2_X1 \mreg/_10506_ ( .A(\mreg/_04417_ ), .B(\mreg/_04966_ ), .S(\mreg/_03830_ ), .Z(\mreg/_00803_ ) );
MUX2_X1 \mreg/_10507_ ( .A(\mreg/_04418_ ), .B(\mreg/_04967_ ), .S(\mreg/_03830_ ), .Z(\mreg/_00804_ ) );
MUX2_X1 \mreg/_10508_ ( .A(\mreg/_04419_ ), .B(\mreg/_04968_ ), .S(\mreg/_03830_ ), .Z(\mreg/_00805_ ) );
MUX2_X1 \mreg/_10509_ ( .A(\mreg/_04420_ ), .B(\mreg/_04969_ ), .S(\mreg/_03830_ ), .Z(\mreg/_00806_ ) );
MUX2_X1 \mreg/_10510_ ( .A(\mreg/_04421_ ), .B(\mreg/_04970_ ), .S(\mreg/_03830_ ), .Z(\mreg/_00807_ ) );
BUF_X4 \mreg/_10511_ ( .A(\mreg/_03829_ ), .Z(\mreg/_03831_ ) );
MUX2_X1 \mreg/_10512_ ( .A(\mreg/_04391_ ), .B(\mreg/_04940_ ), .S(\mreg/_03831_ ), .Z(\mreg/_00808_ ) );
MUX2_X1 \mreg/_10513_ ( .A(\mreg/_04392_ ), .B(\mreg/_04941_ ), .S(\mreg/_03831_ ), .Z(\mreg/_00809_ ) );
MUX2_X1 \mreg/_10514_ ( .A(\mreg/_04393_ ), .B(\mreg/_04942_ ), .S(\mreg/_03831_ ), .Z(\mreg/_00810_ ) );
MUX2_X1 \mreg/_10515_ ( .A(\mreg/_04394_ ), .B(\mreg/_04943_ ), .S(\mreg/_03831_ ), .Z(\mreg/_00811_ ) );
MUX2_X1 \mreg/_10516_ ( .A(\mreg/_04395_ ), .B(\mreg/_04944_ ), .S(\mreg/_03831_ ), .Z(\mreg/_00812_ ) );
MUX2_X1 \mreg/_10517_ ( .A(\mreg/_04396_ ), .B(\mreg/_04945_ ), .S(\mreg/_03831_ ), .Z(\mreg/_00813_ ) );
MUX2_X1 \mreg/_10518_ ( .A(\mreg/_04397_ ), .B(\mreg/_04946_ ), .S(\mreg/_03831_ ), .Z(\mreg/_00814_ ) );
MUX2_X1 \mreg/_10519_ ( .A(\mreg/_04398_ ), .B(\mreg/_04947_ ), .S(\mreg/_03831_ ), .Z(\mreg/_00815_ ) );
MUX2_X1 \mreg/_10520_ ( .A(\mreg/_04399_ ), .B(\mreg/_04948_ ), .S(\mreg/_03831_ ), .Z(\mreg/_00816_ ) );
MUX2_X1 \mreg/_10521_ ( .A(\mreg/_04400_ ), .B(\mreg/_04949_ ), .S(\mreg/_03831_ ), .Z(\mreg/_00817_ ) );
BUF_X4 \mreg/_10522_ ( .A(\mreg/_03829_ ), .Z(\mreg/_03832_ ) );
MUX2_X1 \mreg/_10523_ ( .A(\mreg/_04402_ ), .B(\mreg/_04951_ ), .S(\mreg/_03832_ ), .Z(\mreg/_00818_ ) );
MUX2_X1 \mreg/_10524_ ( .A(\mreg/_04403_ ), .B(\mreg/_04952_ ), .S(\mreg/_03832_ ), .Z(\mreg/_00819_ ) );
MUX2_X1 \mreg/_10525_ ( .A(\mreg/_04404_ ), .B(\mreg/_04953_ ), .S(\mreg/_03832_ ), .Z(\mreg/_00820_ ) );
MUX2_X1 \mreg/_10526_ ( .A(\mreg/_04405_ ), .B(\mreg/_04954_ ), .S(\mreg/_03832_ ), .Z(\mreg/_00821_ ) );
MUX2_X1 \mreg/_10527_ ( .A(\mreg/_04406_ ), .B(\mreg/_04955_ ), .S(\mreg/_03832_ ), .Z(\mreg/_00822_ ) );
MUX2_X1 \mreg/_10528_ ( .A(\mreg/_04407_ ), .B(\mreg/_04956_ ), .S(\mreg/_03832_ ), .Z(\mreg/_00823_ ) );
MUX2_X1 \mreg/_10529_ ( .A(\mreg/_04408_ ), .B(\mreg/_04957_ ), .S(\mreg/_03832_ ), .Z(\mreg/_00824_ ) );
MUX2_X1 \mreg/_10530_ ( .A(\mreg/_04409_ ), .B(\mreg/_04958_ ), .S(\mreg/_03832_ ), .Z(\mreg/_00825_ ) );
MUX2_X1 \mreg/_10531_ ( .A(\mreg/_04410_ ), .B(\mreg/_04959_ ), .S(\mreg/_03832_ ), .Z(\mreg/_00826_ ) );
MUX2_X1 \mreg/_10532_ ( .A(\mreg/_04411_ ), .B(\mreg/_04960_ ), .S(\mreg/_03832_ ), .Z(\mreg/_00827_ ) );
MUX2_X1 \mreg/_10533_ ( .A(\mreg/_04413_ ), .B(\mreg/_04962_ ), .S(\mreg/_03829_ ), .Z(\mreg/_00828_ ) );
MUX2_X1 \mreg/_10534_ ( .A(\mreg/_04414_ ), .B(\mreg/_04963_ ), .S(\mreg/_03829_ ), .Z(\mreg/_00829_ ) );
NAND4_X1 \mreg/_10535_ ( .A1(\mreg/_03691_ ), .A2(\mreg/_04938_ ), .A3(\mreg/_03725_ ), .A4(\mreg/_04937_ ), .ZN(\mreg/_03833_ ) );
NOR2_X1 \mreg/_10536_ ( .A1(\mreg/_03696_ ), .A2(\mreg/_03833_ ), .ZN(\mreg/_03834_ ) );
BUF_X4 \mreg/_10537_ ( .A(\mreg/_03834_ ), .Z(\mreg/_03835_ ) );
MUX2_X1 \mreg/_10538_ ( .A(\mreg/_04422_ ), .B(\mreg/_04939_ ), .S(\mreg/_03835_ ), .Z(\mreg/_00830_ ) );
MUX2_X1 \mreg/_10539_ ( .A(\mreg/_04433_ ), .B(\mreg/_04950_ ), .S(\mreg/_03835_ ), .Z(\mreg/_00831_ ) );
MUX2_X1 \mreg/_10540_ ( .A(\mreg/_04444_ ), .B(\mreg/_04961_ ), .S(\mreg/_03835_ ), .Z(\mreg/_00832_ ) );
MUX2_X1 \mreg/_10541_ ( .A(\mreg/_04447_ ), .B(\mreg/_04964_ ), .S(\mreg/_03835_ ), .Z(\mreg/_00833_ ) );
MUX2_X1 \mreg/_10542_ ( .A(\mreg/_04448_ ), .B(\mreg/_04965_ ), .S(\mreg/_03835_ ), .Z(\mreg/_00834_ ) );
MUX2_X1 \mreg/_10543_ ( .A(\mreg/_04449_ ), .B(\mreg/_04966_ ), .S(\mreg/_03835_ ), .Z(\mreg/_00835_ ) );
MUX2_X1 \mreg/_10544_ ( .A(\mreg/_04450_ ), .B(\mreg/_04967_ ), .S(\mreg/_03835_ ), .Z(\mreg/_00836_ ) );
MUX2_X1 \mreg/_10545_ ( .A(\mreg/_04451_ ), .B(\mreg/_04968_ ), .S(\mreg/_03835_ ), .Z(\mreg/_00837_ ) );
MUX2_X1 \mreg/_10546_ ( .A(\mreg/_04452_ ), .B(\mreg/_04969_ ), .S(\mreg/_03835_ ), .Z(\mreg/_00838_ ) );
MUX2_X1 \mreg/_10547_ ( .A(\mreg/_04453_ ), .B(\mreg/_04970_ ), .S(\mreg/_03835_ ), .Z(\mreg/_00839_ ) );
BUF_X4 \mreg/_10548_ ( .A(\mreg/_03834_ ), .Z(\mreg/_03836_ ) );
MUX2_X1 \mreg/_10549_ ( .A(\mreg/_04423_ ), .B(\mreg/_04940_ ), .S(\mreg/_03836_ ), .Z(\mreg/_00840_ ) );
MUX2_X1 \mreg/_10550_ ( .A(\mreg/_04424_ ), .B(\mreg/_04941_ ), .S(\mreg/_03836_ ), .Z(\mreg/_00841_ ) );
MUX2_X1 \mreg/_10551_ ( .A(\mreg/_04425_ ), .B(\mreg/_04942_ ), .S(\mreg/_03836_ ), .Z(\mreg/_00842_ ) );
MUX2_X1 \mreg/_10552_ ( .A(\mreg/_04426_ ), .B(\mreg/_04943_ ), .S(\mreg/_03836_ ), .Z(\mreg/_00843_ ) );
MUX2_X1 \mreg/_10553_ ( .A(\mreg/_04427_ ), .B(\mreg/_04944_ ), .S(\mreg/_03836_ ), .Z(\mreg/_00844_ ) );
MUX2_X1 \mreg/_10554_ ( .A(\mreg/_04428_ ), .B(\mreg/_04945_ ), .S(\mreg/_03836_ ), .Z(\mreg/_00845_ ) );
MUX2_X1 \mreg/_10555_ ( .A(\mreg/_04429_ ), .B(\mreg/_04946_ ), .S(\mreg/_03836_ ), .Z(\mreg/_00846_ ) );
MUX2_X1 \mreg/_10556_ ( .A(\mreg/_04430_ ), .B(\mreg/_04947_ ), .S(\mreg/_03836_ ), .Z(\mreg/_00847_ ) );
MUX2_X1 \mreg/_10557_ ( .A(\mreg/_04431_ ), .B(\mreg/_04948_ ), .S(\mreg/_03836_ ), .Z(\mreg/_00848_ ) );
MUX2_X1 \mreg/_10558_ ( .A(\mreg/_04432_ ), .B(\mreg/_04949_ ), .S(\mreg/_03836_ ), .Z(\mreg/_00849_ ) );
BUF_X4 \mreg/_10559_ ( .A(\mreg/_03834_ ), .Z(\mreg/_03837_ ) );
MUX2_X1 \mreg/_10560_ ( .A(\mreg/_04434_ ), .B(\mreg/_04951_ ), .S(\mreg/_03837_ ), .Z(\mreg/_00850_ ) );
MUX2_X1 \mreg/_10561_ ( .A(\mreg/_04435_ ), .B(\mreg/_04952_ ), .S(\mreg/_03837_ ), .Z(\mreg/_00851_ ) );
MUX2_X1 \mreg/_10562_ ( .A(\mreg/_04436_ ), .B(\mreg/_04953_ ), .S(\mreg/_03837_ ), .Z(\mreg/_00852_ ) );
MUX2_X1 \mreg/_10563_ ( .A(\mreg/_04437_ ), .B(\mreg/_04954_ ), .S(\mreg/_03837_ ), .Z(\mreg/_00853_ ) );
MUX2_X1 \mreg/_10564_ ( .A(\mreg/_04438_ ), .B(\mreg/_04955_ ), .S(\mreg/_03837_ ), .Z(\mreg/_00854_ ) );
MUX2_X1 \mreg/_10565_ ( .A(\mreg/_04439_ ), .B(\mreg/_04956_ ), .S(\mreg/_03837_ ), .Z(\mreg/_00855_ ) );
MUX2_X1 \mreg/_10566_ ( .A(\mreg/_04440_ ), .B(\mreg/_04957_ ), .S(\mreg/_03837_ ), .Z(\mreg/_00856_ ) );
MUX2_X1 \mreg/_10567_ ( .A(\mreg/_04441_ ), .B(\mreg/_04958_ ), .S(\mreg/_03837_ ), .Z(\mreg/_00857_ ) );
MUX2_X1 \mreg/_10568_ ( .A(\mreg/_04442_ ), .B(\mreg/_04959_ ), .S(\mreg/_03837_ ), .Z(\mreg/_00858_ ) );
MUX2_X1 \mreg/_10569_ ( .A(\mreg/_04443_ ), .B(\mreg/_04960_ ), .S(\mreg/_03837_ ), .Z(\mreg/_00859_ ) );
MUX2_X1 \mreg/_10570_ ( .A(\mreg/_04445_ ), .B(\mreg/_04962_ ), .S(\mreg/_03834_ ), .Z(\mreg/_00860_ ) );
MUX2_X1 \mreg/_10571_ ( .A(\mreg/_04446_ ), .B(\mreg/_04963_ ), .S(\mreg/_03834_ ), .Z(\mreg/_00861_ ) );
OR3_X1 \mreg/_10572_ ( .A1(\mreg/_03706_ ), .A2(\mreg/_03714_ ), .A3(\mreg/_03755_ ), .ZN(\mreg/_03838_ ) );
NOR2_X1 \mreg/_10573_ ( .A1(\mreg/_03838_ ), .A2(\mreg/_03783_ ), .ZN(\mreg/_03839_ ) );
BUF_X4 \mreg/_10574_ ( .A(\mreg/_03839_ ), .Z(\mreg/_03840_ ) );
MUX2_X1 \mreg/_10575_ ( .A(\mreg/_04454_ ), .B(\mreg/_04939_ ), .S(\mreg/_03840_ ), .Z(\mreg/_00862_ ) );
MUX2_X1 \mreg/_10576_ ( .A(\mreg/_04465_ ), .B(\mreg/_04950_ ), .S(\mreg/_03840_ ), .Z(\mreg/_00863_ ) );
MUX2_X1 \mreg/_10577_ ( .A(\mreg/_04476_ ), .B(\mreg/_04961_ ), .S(\mreg/_03840_ ), .Z(\mreg/_00864_ ) );
MUX2_X1 \mreg/_10578_ ( .A(\mreg/_04479_ ), .B(\mreg/_04964_ ), .S(\mreg/_03840_ ), .Z(\mreg/_00865_ ) );
MUX2_X1 \mreg/_10579_ ( .A(\mreg/_04480_ ), .B(\mreg/_04965_ ), .S(\mreg/_03840_ ), .Z(\mreg/_00866_ ) );
MUX2_X1 \mreg/_10580_ ( .A(\mreg/_04481_ ), .B(\mreg/_04966_ ), .S(\mreg/_03840_ ), .Z(\mreg/_00867_ ) );
MUX2_X1 \mreg/_10581_ ( .A(\mreg/_04482_ ), .B(\mreg/_04967_ ), .S(\mreg/_03840_ ), .Z(\mreg/_00868_ ) );
MUX2_X1 \mreg/_10582_ ( .A(\mreg/_04483_ ), .B(\mreg/_04968_ ), .S(\mreg/_03840_ ), .Z(\mreg/_00869_ ) );
MUX2_X1 \mreg/_10583_ ( .A(\mreg/_04484_ ), .B(\mreg/_04969_ ), .S(\mreg/_03840_ ), .Z(\mreg/_00870_ ) );
MUX2_X1 \mreg/_10584_ ( .A(\mreg/_04485_ ), .B(\mreg/_04970_ ), .S(\mreg/_03840_ ), .Z(\mreg/_00871_ ) );
BUF_X4 \mreg/_10585_ ( .A(\mreg/_03839_ ), .Z(\mreg/_03841_ ) );
MUX2_X1 \mreg/_10586_ ( .A(\mreg/_04455_ ), .B(\mreg/_04940_ ), .S(\mreg/_03841_ ), .Z(\mreg/_00872_ ) );
MUX2_X1 \mreg/_10587_ ( .A(\mreg/_04456_ ), .B(\mreg/_04941_ ), .S(\mreg/_03841_ ), .Z(\mreg/_00873_ ) );
MUX2_X1 \mreg/_10588_ ( .A(\mreg/_04457_ ), .B(\mreg/_04942_ ), .S(\mreg/_03841_ ), .Z(\mreg/_00874_ ) );
MUX2_X1 \mreg/_10589_ ( .A(\mreg/_04458_ ), .B(\mreg/_04943_ ), .S(\mreg/_03841_ ), .Z(\mreg/_00875_ ) );
MUX2_X1 \mreg/_10590_ ( .A(\mreg/_04459_ ), .B(\mreg/_04944_ ), .S(\mreg/_03841_ ), .Z(\mreg/_00876_ ) );
MUX2_X1 \mreg/_10591_ ( .A(\mreg/_04460_ ), .B(\mreg/_04945_ ), .S(\mreg/_03841_ ), .Z(\mreg/_00877_ ) );
MUX2_X1 \mreg/_10592_ ( .A(\mreg/_04461_ ), .B(\mreg/_04946_ ), .S(\mreg/_03841_ ), .Z(\mreg/_00878_ ) );
MUX2_X1 \mreg/_10593_ ( .A(\mreg/_04462_ ), .B(\mreg/_04947_ ), .S(\mreg/_03841_ ), .Z(\mreg/_00879_ ) );
MUX2_X1 \mreg/_10594_ ( .A(\mreg/_04463_ ), .B(\mreg/_04948_ ), .S(\mreg/_03841_ ), .Z(\mreg/_00880_ ) );
MUX2_X1 \mreg/_10595_ ( .A(\mreg/_04464_ ), .B(\mreg/_04949_ ), .S(\mreg/_03841_ ), .Z(\mreg/_00881_ ) );
BUF_X4 \mreg/_10596_ ( .A(\mreg/_03839_ ), .Z(\mreg/_03842_ ) );
MUX2_X1 \mreg/_10597_ ( .A(\mreg/_04466_ ), .B(\mreg/_04951_ ), .S(\mreg/_03842_ ), .Z(\mreg/_00882_ ) );
MUX2_X1 \mreg/_10598_ ( .A(\mreg/_04467_ ), .B(\mreg/_04952_ ), .S(\mreg/_03842_ ), .Z(\mreg/_00883_ ) );
MUX2_X1 \mreg/_10599_ ( .A(\mreg/_04468_ ), .B(\mreg/_04953_ ), .S(\mreg/_03842_ ), .Z(\mreg/_00884_ ) );
MUX2_X1 \mreg/_10600_ ( .A(\mreg/_04469_ ), .B(\mreg/_04954_ ), .S(\mreg/_03842_ ), .Z(\mreg/_00885_ ) );
MUX2_X1 \mreg/_10601_ ( .A(\mreg/_04470_ ), .B(\mreg/_04955_ ), .S(\mreg/_03842_ ), .Z(\mreg/_00886_ ) );
MUX2_X1 \mreg/_10602_ ( .A(\mreg/_04471_ ), .B(\mreg/_04956_ ), .S(\mreg/_03842_ ), .Z(\mreg/_00887_ ) );
MUX2_X1 \mreg/_10603_ ( .A(\mreg/_04472_ ), .B(\mreg/_04957_ ), .S(\mreg/_03842_ ), .Z(\mreg/_00888_ ) );
MUX2_X1 \mreg/_10604_ ( .A(\mreg/_04473_ ), .B(\mreg/_04958_ ), .S(\mreg/_03842_ ), .Z(\mreg/_00889_ ) );
MUX2_X1 \mreg/_10605_ ( .A(\mreg/_04474_ ), .B(\mreg/_04959_ ), .S(\mreg/_03842_ ), .Z(\mreg/_00890_ ) );
MUX2_X1 \mreg/_10606_ ( .A(\mreg/_04475_ ), .B(\mreg/_04960_ ), .S(\mreg/_03842_ ), .Z(\mreg/_00891_ ) );
MUX2_X1 \mreg/_10607_ ( .A(\mreg/_04477_ ), .B(\mreg/_04962_ ), .S(\mreg/_03839_ ), .Z(\mreg/_00892_ ) );
MUX2_X1 \mreg/_10608_ ( .A(\mreg/_04478_ ), .B(\mreg/_04963_ ), .S(\mreg/_03839_ ), .Z(\mreg/_00893_ ) );
NAND2_X1 \mreg/_10609_ ( .A1(\mreg/_03761_ ), .A2(\mreg/_04938_ ), .ZN(\mreg/_03843_ ) );
NOR2_X1 \mreg/_10610_ ( .A1(\mreg/_03843_ ), .A2(\mreg/_03783_ ), .ZN(\mreg/_03844_ ) );
BUF_X4 \mreg/_10611_ ( .A(\mreg/_03844_ ), .Z(\mreg/_03845_ ) );
MUX2_X1 \mreg/_10612_ ( .A(\mreg/_04486_ ), .B(\mreg/_04939_ ), .S(\mreg/_03845_ ), .Z(\mreg/_00894_ ) );
MUX2_X1 \mreg/_10613_ ( .A(\mreg/_04497_ ), .B(\mreg/_04950_ ), .S(\mreg/_03845_ ), .Z(\mreg/_00895_ ) );
MUX2_X1 \mreg/_10614_ ( .A(\mreg/_04508_ ), .B(\mreg/_04961_ ), .S(\mreg/_03845_ ), .Z(\mreg/_00896_ ) );
MUX2_X1 \mreg/_10615_ ( .A(\mreg/_04511_ ), .B(\mreg/_04964_ ), .S(\mreg/_03845_ ), .Z(\mreg/_00897_ ) );
MUX2_X1 \mreg/_10616_ ( .A(\mreg/_04512_ ), .B(\mreg/_04965_ ), .S(\mreg/_03845_ ), .Z(\mreg/_00898_ ) );
MUX2_X1 \mreg/_10617_ ( .A(\mreg/_04513_ ), .B(\mreg/_04966_ ), .S(\mreg/_03845_ ), .Z(\mreg/_00899_ ) );
MUX2_X1 \mreg/_10618_ ( .A(\mreg/_04514_ ), .B(\mreg/_04967_ ), .S(\mreg/_03845_ ), .Z(\mreg/_00900_ ) );
MUX2_X1 \mreg/_10619_ ( .A(\mreg/_04515_ ), .B(\mreg/_04968_ ), .S(\mreg/_03845_ ), .Z(\mreg/_00901_ ) );
MUX2_X1 \mreg/_10620_ ( .A(\mreg/_04516_ ), .B(\mreg/_04969_ ), .S(\mreg/_03845_ ), .Z(\mreg/_00902_ ) );
MUX2_X1 \mreg/_10621_ ( .A(\mreg/_04517_ ), .B(\mreg/_04970_ ), .S(\mreg/_03845_ ), .Z(\mreg/_00903_ ) );
BUF_X4 \mreg/_10622_ ( .A(\mreg/_03844_ ), .Z(\mreg/_03846_ ) );
MUX2_X1 \mreg/_10623_ ( .A(\mreg/_04487_ ), .B(\mreg/_04940_ ), .S(\mreg/_03846_ ), .Z(\mreg/_00904_ ) );
MUX2_X1 \mreg/_10624_ ( .A(\mreg/_04488_ ), .B(\mreg/_04941_ ), .S(\mreg/_03846_ ), .Z(\mreg/_00905_ ) );
MUX2_X1 \mreg/_10625_ ( .A(\mreg/_04489_ ), .B(\mreg/_04942_ ), .S(\mreg/_03846_ ), .Z(\mreg/_00906_ ) );
MUX2_X1 \mreg/_10626_ ( .A(\mreg/_04490_ ), .B(\mreg/_04943_ ), .S(\mreg/_03846_ ), .Z(\mreg/_00907_ ) );
MUX2_X1 \mreg/_10627_ ( .A(\mreg/_04491_ ), .B(\mreg/_04944_ ), .S(\mreg/_03846_ ), .Z(\mreg/_00908_ ) );
MUX2_X1 \mreg/_10628_ ( .A(\mreg/_04492_ ), .B(\mreg/_04945_ ), .S(\mreg/_03846_ ), .Z(\mreg/_00909_ ) );
MUX2_X1 \mreg/_10629_ ( .A(\mreg/_04493_ ), .B(\mreg/_04946_ ), .S(\mreg/_03846_ ), .Z(\mreg/_00910_ ) );
MUX2_X1 \mreg/_10630_ ( .A(\mreg/_04494_ ), .B(\mreg/_04947_ ), .S(\mreg/_03846_ ), .Z(\mreg/_00911_ ) );
MUX2_X1 \mreg/_10631_ ( .A(\mreg/_04495_ ), .B(\mreg/_04948_ ), .S(\mreg/_03846_ ), .Z(\mreg/_00912_ ) );
MUX2_X1 \mreg/_10632_ ( .A(\mreg/_04496_ ), .B(\mreg/_04949_ ), .S(\mreg/_03846_ ), .Z(\mreg/_00913_ ) );
BUF_X4 \mreg/_10633_ ( .A(\mreg/_03844_ ), .Z(\mreg/_03847_ ) );
MUX2_X1 \mreg/_10634_ ( .A(\mreg/_04498_ ), .B(\mreg/_04951_ ), .S(\mreg/_03847_ ), .Z(\mreg/_00914_ ) );
MUX2_X1 \mreg/_10635_ ( .A(\mreg/_04499_ ), .B(\mreg/_04952_ ), .S(\mreg/_03847_ ), .Z(\mreg/_00915_ ) );
MUX2_X1 \mreg/_10636_ ( .A(\mreg/_04500_ ), .B(\mreg/_04953_ ), .S(\mreg/_03847_ ), .Z(\mreg/_00916_ ) );
MUX2_X1 \mreg/_10637_ ( .A(\mreg/_04501_ ), .B(\mreg/_04954_ ), .S(\mreg/_03847_ ), .Z(\mreg/_00917_ ) );
MUX2_X1 \mreg/_10638_ ( .A(\mreg/_04502_ ), .B(\mreg/_04955_ ), .S(\mreg/_03847_ ), .Z(\mreg/_00918_ ) );
MUX2_X1 \mreg/_10639_ ( .A(\mreg/_04503_ ), .B(\mreg/_04956_ ), .S(\mreg/_03847_ ), .Z(\mreg/_00919_ ) );
MUX2_X1 \mreg/_10640_ ( .A(\mreg/_04504_ ), .B(\mreg/_04957_ ), .S(\mreg/_03847_ ), .Z(\mreg/_00920_ ) );
MUX2_X1 \mreg/_10641_ ( .A(\mreg/_04505_ ), .B(\mreg/_04958_ ), .S(\mreg/_03847_ ), .Z(\mreg/_00921_ ) );
MUX2_X1 \mreg/_10642_ ( .A(\mreg/_04506_ ), .B(\mreg/_04959_ ), .S(\mreg/_03847_ ), .Z(\mreg/_00922_ ) );
MUX2_X1 \mreg/_10643_ ( .A(\mreg/_04507_ ), .B(\mreg/_04960_ ), .S(\mreg/_03847_ ), .Z(\mreg/_00923_ ) );
MUX2_X1 \mreg/_10644_ ( .A(\mreg/_04509_ ), .B(\mreg/_04962_ ), .S(\mreg/_03844_ ), .Z(\mreg/_00924_ ) );
MUX2_X1 \mreg/_10645_ ( .A(\mreg/_04510_ ), .B(\mreg/_04963_ ), .S(\mreg/_03844_ ), .Z(\mreg/_00925_ ) );
OR3_X1 \mreg/_10646_ ( .A1(\mreg/_03755_ ), .A2(\mreg/_03714_ ), .A3(\mreg/_03698_ ), .ZN(\mreg/_03848_ ) );
NOR2_X1 \mreg/_10647_ ( .A1(\mreg/_03848_ ), .A2(\mreg/_03783_ ), .ZN(\mreg/_03849_ ) );
BUF_X4 \mreg/_10648_ ( .A(\mreg/_03849_ ), .Z(\mreg/_03850_ ) );
MUX2_X1 \mreg/_10649_ ( .A(\mreg/_04518_ ), .B(\mreg/_04939_ ), .S(\mreg/_03850_ ), .Z(\mreg/_00926_ ) );
MUX2_X1 \mreg/_10650_ ( .A(\mreg/_04529_ ), .B(\mreg/_04950_ ), .S(\mreg/_03850_ ), .Z(\mreg/_00927_ ) );
MUX2_X1 \mreg/_10651_ ( .A(\mreg/_04540_ ), .B(\mreg/_04961_ ), .S(\mreg/_03850_ ), .Z(\mreg/_00928_ ) );
MUX2_X1 \mreg/_10652_ ( .A(\mreg/_04543_ ), .B(\mreg/_04964_ ), .S(\mreg/_03850_ ), .Z(\mreg/_00929_ ) );
MUX2_X1 \mreg/_10653_ ( .A(\mreg/_04544_ ), .B(\mreg/_04965_ ), .S(\mreg/_03850_ ), .Z(\mreg/_00930_ ) );
MUX2_X1 \mreg/_10654_ ( .A(\mreg/_04545_ ), .B(\mreg/_04966_ ), .S(\mreg/_03850_ ), .Z(\mreg/_00931_ ) );
MUX2_X1 \mreg/_10655_ ( .A(\mreg/_04546_ ), .B(\mreg/_04967_ ), .S(\mreg/_03850_ ), .Z(\mreg/_00932_ ) );
MUX2_X1 \mreg/_10656_ ( .A(\mreg/_04547_ ), .B(\mreg/_04968_ ), .S(\mreg/_03850_ ), .Z(\mreg/_00933_ ) );
MUX2_X1 \mreg/_10657_ ( .A(\mreg/_04548_ ), .B(\mreg/_04969_ ), .S(\mreg/_03850_ ), .Z(\mreg/_00934_ ) );
MUX2_X1 \mreg/_10658_ ( .A(\mreg/_04549_ ), .B(\mreg/_04970_ ), .S(\mreg/_03850_ ), .Z(\mreg/_00935_ ) );
BUF_X4 \mreg/_10659_ ( .A(\mreg/_03849_ ), .Z(\mreg/_03851_ ) );
MUX2_X1 \mreg/_10660_ ( .A(\mreg/_04519_ ), .B(\mreg/_04940_ ), .S(\mreg/_03851_ ), .Z(\mreg/_00936_ ) );
MUX2_X1 \mreg/_10661_ ( .A(\mreg/_04520_ ), .B(\mreg/_04941_ ), .S(\mreg/_03851_ ), .Z(\mreg/_00937_ ) );
MUX2_X1 \mreg/_10662_ ( .A(\mreg/_04521_ ), .B(\mreg/_04942_ ), .S(\mreg/_03851_ ), .Z(\mreg/_00938_ ) );
MUX2_X1 \mreg/_10663_ ( .A(\mreg/_04522_ ), .B(\mreg/_04943_ ), .S(\mreg/_03851_ ), .Z(\mreg/_00939_ ) );
MUX2_X1 \mreg/_10664_ ( .A(\mreg/_04523_ ), .B(\mreg/_04944_ ), .S(\mreg/_03851_ ), .Z(\mreg/_00940_ ) );
MUX2_X1 \mreg/_10665_ ( .A(\mreg/_04524_ ), .B(\mreg/_04945_ ), .S(\mreg/_03851_ ), .Z(\mreg/_00941_ ) );
MUX2_X1 \mreg/_10666_ ( .A(\mreg/_04525_ ), .B(\mreg/_04946_ ), .S(\mreg/_03851_ ), .Z(\mreg/_00942_ ) );
MUX2_X1 \mreg/_10667_ ( .A(\mreg/_04526_ ), .B(\mreg/_04947_ ), .S(\mreg/_03851_ ), .Z(\mreg/_00943_ ) );
MUX2_X1 \mreg/_10668_ ( .A(\mreg/_04527_ ), .B(\mreg/_04948_ ), .S(\mreg/_03851_ ), .Z(\mreg/_00944_ ) );
MUX2_X1 \mreg/_10669_ ( .A(\mreg/_04528_ ), .B(\mreg/_04949_ ), .S(\mreg/_03851_ ), .Z(\mreg/_00945_ ) );
BUF_X4 \mreg/_10670_ ( .A(\mreg/_03849_ ), .Z(\mreg/_03852_ ) );
MUX2_X1 \mreg/_10671_ ( .A(\mreg/_04530_ ), .B(\mreg/_04951_ ), .S(\mreg/_03852_ ), .Z(\mreg/_00946_ ) );
MUX2_X1 \mreg/_10672_ ( .A(\mreg/_04531_ ), .B(\mreg/_04952_ ), .S(\mreg/_03852_ ), .Z(\mreg/_00947_ ) );
MUX2_X1 \mreg/_10673_ ( .A(\mreg/_04532_ ), .B(\mreg/_04953_ ), .S(\mreg/_03852_ ), .Z(\mreg/_00948_ ) );
MUX2_X1 \mreg/_10674_ ( .A(\mreg/_04533_ ), .B(\mreg/_04954_ ), .S(\mreg/_03852_ ), .Z(\mreg/_00949_ ) );
MUX2_X1 \mreg/_10675_ ( .A(\mreg/_04534_ ), .B(\mreg/_04955_ ), .S(\mreg/_03852_ ), .Z(\mreg/_00950_ ) );
MUX2_X1 \mreg/_10676_ ( .A(\mreg/_04535_ ), .B(\mreg/_04956_ ), .S(\mreg/_03852_ ), .Z(\mreg/_00951_ ) );
MUX2_X1 \mreg/_10677_ ( .A(\mreg/_04536_ ), .B(\mreg/_04957_ ), .S(\mreg/_03852_ ), .Z(\mreg/_00952_ ) );
MUX2_X1 \mreg/_10678_ ( .A(\mreg/_04537_ ), .B(\mreg/_04958_ ), .S(\mreg/_03852_ ), .Z(\mreg/_00953_ ) );
MUX2_X1 \mreg/_10679_ ( .A(\mreg/_04538_ ), .B(\mreg/_04959_ ), .S(\mreg/_03852_ ), .Z(\mreg/_00954_ ) );
MUX2_X1 \mreg/_10680_ ( .A(\mreg/_04539_ ), .B(\mreg/_04960_ ), .S(\mreg/_03852_ ), .Z(\mreg/_00955_ ) );
MUX2_X1 \mreg/_10681_ ( .A(\mreg/_04541_ ), .B(\mreg/_04962_ ), .S(\mreg/_03849_ ), .Z(\mreg/_00956_ ) );
MUX2_X1 \mreg/_10682_ ( .A(\mreg/_04542_ ), .B(\mreg/_04963_ ), .S(\mreg/_03849_ ), .Z(\mreg/_00957_ ) );
NAND4_X1 \mreg/_10683_ ( .A1(\mreg/_03691_ ), .A2(\mreg/_04938_ ), .A3(\mreg/_04936_ ), .A4(\mreg/_04937_ ), .ZN(\mreg/_03853_ ) );
NOR2_X1 \mreg/_10684_ ( .A1(\mreg/_03709_ ), .A2(\mreg/_03853_ ), .ZN(\mreg/_03854_ ) );
BUF_X4 \mreg/_10685_ ( .A(\mreg/_03854_ ), .Z(\mreg/_03855_ ) );
MUX2_X1 \mreg/_10686_ ( .A(\mreg/_04550_ ), .B(\mreg/_04939_ ), .S(\mreg/_03855_ ), .Z(\mreg/_00958_ ) );
MUX2_X1 \mreg/_10687_ ( .A(\mreg/_04561_ ), .B(\mreg/_04950_ ), .S(\mreg/_03855_ ), .Z(\mreg/_00959_ ) );
MUX2_X1 \mreg/_10688_ ( .A(\mreg/_04572_ ), .B(\mreg/_04961_ ), .S(\mreg/_03855_ ), .Z(\mreg/_00960_ ) );
MUX2_X1 \mreg/_10689_ ( .A(\mreg/_04575_ ), .B(\mreg/_04964_ ), .S(\mreg/_03855_ ), .Z(\mreg/_00961_ ) );
MUX2_X1 \mreg/_10690_ ( .A(\mreg/_04576_ ), .B(\mreg/_04965_ ), .S(\mreg/_03855_ ), .Z(\mreg/_00962_ ) );
MUX2_X1 \mreg/_10691_ ( .A(\mreg/_04577_ ), .B(\mreg/_04966_ ), .S(\mreg/_03855_ ), .Z(\mreg/_00963_ ) );
MUX2_X1 \mreg/_10692_ ( .A(\mreg/_04578_ ), .B(\mreg/_04967_ ), .S(\mreg/_03855_ ), .Z(\mreg/_00964_ ) );
MUX2_X1 \mreg/_10693_ ( .A(\mreg/_04579_ ), .B(\mreg/_04968_ ), .S(\mreg/_03855_ ), .Z(\mreg/_00965_ ) );
MUX2_X1 \mreg/_10694_ ( .A(\mreg/_04580_ ), .B(\mreg/_04969_ ), .S(\mreg/_03855_ ), .Z(\mreg/_00966_ ) );
MUX2_X1 \mreg/_10695_ ( .A(\mreg/_04581_ ), .B(\mreg/_04970_ ), .S(\mreg/_03855_ ), .Z(\mreg/_00967_ ) );
BUF_X4 \mreg/_10696_ ( .A(\mreg/_03854_ ), .Z(\mreg/_03856_ ) );
MUX2_X1 \mreg/_10697_ ( .A(\mreg/_04551_ ), .B(\mreg/_04940_ ), .S(\mreg/_03856_ ), .Z(\mreg/_00968_ ) );
MUX2_X1 \mreg/_10698_ ( .A(\mreg/_04552_ ), .B(\mreg/_04941_ ), .S(\mreg/_03856_ ), .Z(\mreg/_00969_ ) );
MUX2_X1 \mreg/_10699_ ( .A(\mreg/_04553_ ), .B(\mreg/_04942_ ), .S(\mreg/_03856_ ), .Z(\mreg/_00970_ ) );
MUX2_X1 \mreg/_10700_ ( .A(\mreg/_04554_ ), .B(\mreg/_04943_ ), .S(\mreg/_03856_ ), .Z(\mreg/_00971_ ) );
MUX2_X1 \mreg/_10701_ ( .A(\mreg/_04555_ ), .B(\mreg/_04944_ ), .S(\mreg/_03856_ ), .Z(\mreg/_00972_ ) );
MUX2_X1 \mreg/_10702_ ( .A(\mreg/_04556_ ), .B(\mreg/_04945_ ), .S(\mreg/_03856_ ), .Z(\mreg/_00973_ ) );
MUX2_X1 \mreg/_10703_ ( .A(\mreg/_04557_ ), .B(\mreg/_04946_ ), .S(\mreg/_03856_ ), .Z(\mreg/_00974_ ) );
MUX2_X1 \mreg/_10704_ ( .A(\mreg/_04558_ ), .B(\mreg/_04947_ ), .S(\mreg/_03856_ ), .Z(\mreg/_00975_ ) );
MUX2_X1 \mreg/_10705_ ( .A(\mreg/_04559_ ), .B(\mreg/_04948_ ), .S(\mreg/_03856_ ), .Z(\mreg/_00976_ ) );
MUX2_X1 \mreg/_10706_ ( .A(\mreg/_04560_ ), .B(\mreg/_04949_ ), .S(\mreg/_03856_ ), .Z(\mreg/_00977_ ) );
BUF_X4 \mreg/_10707_ ( .A(\mreg/_03854_ ), .Z(\mreg/_03857_ ) );
MUX2_X1 \mreg/_10708_ ( .A(\mreg/_04562_ ), .B(\mreg/_04951_ ), .S(\mreg/_03857_ ), .Z(\mreg/_00978_ ) );
MUX2_X1 \mreg/_10709_ ( .A(\mreg/_04563_ ), .B(\mreg/_04952_ ), .S(\mreg/_03857_ ), .Z(\mreg/_00979_ ) );
MUX2_X1 \mreg/_10710_ ( .A(\mreg/_04564_ ), .B(\mreg/_04953_ ), .S(\mreg/_03857_ ), .Z(\mreg/_00980_ ) );
MUX2_X1 \mreg/_10711_ ( .A(\mreg/_04565_ ), .B(\mreg/_04954_ ), .S(\mreg/_03857_ ), .Z(\mreg/_00981_ ) );
MUX2_X1 \mreg/_10712_ ( .A(\mreg/_04566_ ), .B(\mreg/_04955_ ), .S(\mreg/_03857_ ), .Z(\mreg/_00982_ ) );
MUX2_X1 \mreg/_10713_ ( .A(\mreg/_04567_ ), .B(\mreg/_04956_ ), .S(\mreg/_03857_ ), .Z(\mreg/_00983_ ) );
MUX2_X1 \mreg/_10714_ ( .A(\mreg/_04568_ ), .B(\mreg/_04957_ ), .S(\mreg/_03857_ ), .Z(\mreg/_00984_ ) );
MUX2_X1 \mreg/_10715_ ( .A(\mreg/_04569_ ), .B(\mreg/_04958_ ), .S(\mreg/_03857_ ), .Z(\mreg/_00985_ ) );
MUX2_X1 \mreg/_10716_ ( .A(\mreg/_04570_ ), .B(\mreg/_04959_ ), .S(\mreg/_03857_ ), .Z(\mreg/_00986_ ) );
MUX2_X1 \mreg/_10717_ ( .A(\mreg/_04571_ ), .B(\mreg/_04960_ ), .S(\mreg/_03857_ ), .Z(\mreg/_00987_ ) );
MUX2_X1 \mreg/_10718_ ( .A(\mreg/_04573_ ), .B(\mreg/_04962_ ), .S(\mreg/_03854_ ), .Z(\mreg/_00988_ ) );
MUX2_X1 \mreg/_10719_ ( .A(\mreg/_04574_ ), .B(\mreg/_04963_ ), .S(\mreg/_03854_ ), .Z(\mreg/_00989_ ) );
OR4_X1 \mreg/_10720_ ( .A1(\mreg/_03692_ ), .A2(\mreg/_03697_ ), .A3(\mreg/_03705_ ), .A4(\mreg/_04935_ ), .ZN(\mreg/_03858_ ) );
NOR2_X1 \mreg/_10721_ ( .A1(\mreg/_03858_ ), .A2(\mreg/_03783_ ), .ZN(\mreg/_03859_ ) );
BUF_X4 \mreg/_10722_ ( .A(\mreg/_03859_ ), .Z(\mreg/_03860_ ) );
MUX2_X1 \mreg/_10723_ ( .A(\mreg/_04582_ ), .B(\mreg/_04939_ ), .S(\mreg/_03860_ ), .Z(\mreg/_00990_ ) );
MUX2_X1 \mreg/_10724_ ( .A(\mreg/_04593_ ), .B(\mreg/_04950_ ), .S(\mreg/_03860_ ), .Z(\mreg/_00991_ ) );
MUX2_X1 \mreg/_10725_ ( .A(\mreg/_04604_ ), .B(\mreg/_04961_ ), .S(\mreg/_03860_ ), .Z(\mreg/_00992_ ) );
MUX2_X1 \mreg/_10726_ ( .A(\mreg/_04607_ ), .B(\mreg/_04964_ ), .S(\mreg/_03860_ ), .Z(\mreg/_00993_ ) );
MUX2_X1 \mreg/_10727_ ( .A(\mreg/_04608_ ), .B(\mreg/_04965_ ), .S(\mreg/_03860_ ), .Z(\mreg/_00994_ ) );
MUX2_X1 \mreg/_10728_ ( .A(\mreg/_04609_ ), .B(\mreg/_04966_ ), .S(\mreg/_03860_ ), .Z(\mreg/_00995_ ) );
MUX2_X1 \mreg/_10729_ ( .A(\mreg/_04610_ ), .B(\mreg/_04967_ ), .S(\mreg/_03860_ ), .Z(\mreg/_00996_ ) );
MUX2_X1 \mreg/_10730_ ( .A(\mreg/_04611_ ), .B(\mreg/_04968_ ), .S(\mreg/_03860_ ), .Z(\mreg/_00997_ ) );
MUX2_X1 \mreg/_10731_ ( .A(\mreg/_04612_ ), .B(\mreg/_04969_ ), .S(\mreg/_03860_ ), .Z(\mreg/_00998_ ) );
MUX2_X1 \mreg/_10732_ ( .A(\mreg/_04613_ ), .B(\mreg/_04970_ ), .S(\mreg/_03860_ ), .Z(\mreg/_00999_ ) );
BUF_X4 \mreg/_10733_ ( .A(\mreg/_03859_ ), .Z(\mreg/_03861_ ) );
MUX2_X1 \mreg/_10734_ ( .A(\mreg/_04583_ ), .B(\mreg/_04940_ ), .S(\mreg/_03861_ ), .Z(\mreg/_01000_ ) );
MUX2_X1 \mreg/_10735_ ( .A(\mreg/_04584_ ), .B(\mreg/_04941_ ), .S(\mreg/_03861_ ), .Z(\mreg/_01001_ ) );
MUX2_X1 \mreg/_10736_ ( .A(\mreg/_04585_ ), .B(\mreg/_04942_ ), .S(\mreg/_03861_ ), .Z(\mreg/_01002_ ) );
MUX2_X1 \mreg/_10737_ ( .A(\mreg/_04586_ ), .B(\mreg/_04943_ ), .S(\mreg/_03861_ ), .Z(\mreg/_01003_ ) );
MUX2_X1 \mreg/_10738_ ( .A(\mreg/_04587_ ), .B(\mreg/_04944_ ), .S(\mreg/_03861_ ), .Z(\mreg/_01004_ ) );
MUX2_X1 \mreg/_10739_ ( .A(\mreg/_04588_ ), .B(\mreg/_04945_ ), .S(\mreg/_03861_ ), .Z(\mreg/_01005_ ) );
MUX2_X1 \mreg/_10740_ ( .A(\mreg/_04589_ ), .B(\mreg/_04946_ ), .S(\mreg/_03861_ ), .Z(\mreg/_01006_ ) );
MUX2_X1 \mreg/_10741_ ( .A(\mreg/_04590_ ), .B(\mreg/_04947_ ), .S(\mreg/_03861_ ), .Z(\mreg/_01007_ ) );
MUX2_X1 \mreg/_10742_ ( .A(\mreg/_04591_ ), .B(\mreg/_04948_ ), .S(\mreg/_03861_ ), .Z(\mreg/_01008_ ) );
MUX2_X1 \mreg/_10743_ ( .A(\mreg/_04592_ ), .B(\mreg/_04949_ ), .S(\mreg/_03861_ ), .Z(\mreg/_01009_ ) );
BUF_X4 \mreg/_10744_ ( .A(\mreg/_03859_ ), .Z(\mreg/_03862_ ) );
MUX2_X1 \mreg/_10745_ ( .A(\mreg/_04594_ ), .B(\mreg/_04951_ ), .S(\mreg/_03862_ ), .Z(\mreg/_01010_ ) );
MUX2_X1 \mreg/_10746_ ( .A(\mreg/_04595_ ), .B(\mreg/_04952_ ), .S(\mreg/_03862_ ), .Z(\mreg/_01011_ ) );
MUX2_X1 \mreg/_10747_ ( .A(\mreg/_04596_ ), .B(\mreg/_04953_ ), .S(\mreg/_03862_ ), .Z(\mreg/_01012_ ) );
MUX2_X1 \mreg/_10748_ ( .A(\mreg/_04597_ ), .B(\mreg/_04954_ ), .S(\mreg/_03862_ ), .Z(\mreg/_01013_ ) );
MUX2_X1 \mreg/_10749_ ( .A(\mreg/_04598_ ), .B(\mreg/_04955_ ), .S(\mreg/_03862_ ), .Z(\mreg/_01014_ ) );
MUX2_X1 \mreg/_10750_ ( .A(\mreg/_04599_ ), .B(\mreg/_04956_ ), .S(\mreg/_03862_ ), .Z(\mreg/_01015_ ) );
MUX2_X1 \mreg/_10751_ ( .A(\mreg/_04600_ ), .B(\mreg/_04957_ ), .S(\mreg/_03862_ ), .Z(\mreg/_01016_ ) );
MUX2_X1 \mreg/_10752_ ( .A(\mreg/_04601_ ), .B(\mreg/_04958_ ), .S(\mreg/_03862_ ), .Z(\mreg/_01017_ ) );
MUX2_X1 \mreg/_10753_ ( .A(\mreg/_04602_ ), .B(\mreg/_04959_ ), .S(\mreg/_03862_ ), .Z(\mreg/_01018_ ) );
MUX2_X1 \mreg/_10754_ ( .A(\mreg/_04603_ ), .B(\mreg/_04960_ ), .S(\mreg/_03862_ ), .Z(\mreg/_01019_ ) );
MUX2_X1 \mreg/_10755_ ( .A(\mreg/_04605_ ), .B(\mreg/_04962_ ), .S(\mreg/_03859_ ), .Z(\mreg/_01020_ ) );
MUX2_X1 \mreg/_10756_ ( .A(\mreg/_04606_ ), .B(\mreg/_04963_ ), .S(\mreg/_03859_ ), .Z(\mreg/_01021_ ) );
OR3_X1 \mreg/_10757_ ( .A1(\mreg/_03739_ ), .A2(\mreg/_03692_ ), .A3(\mreg/_03697_ ), .ZN(\mreg/_03863_ ) );
NOR2_X1 \mreg/_10758_ ( .A1(\mreg/_03863_ ), .A2(\mreg/_03695_ ), .ZN(\mreg/_03864_ ) );
BUF_X4 \mreg/_10759_ ( .A(\mreg/_03864_ ), .Z(\mreg/_03865_ ) );
MUX2_X1 \mreg/_10760_ ( .A(\mreg/_04646_ ), .B(\mreg/_04939_ ), .S(\mreg/_03865_ ), .Z(\mreg/_01022_ ) );
MUX2_X1 \mreg/_10761_ ( .A(\mreg/_04657_ ), .B(\mreg/_04950_ ), .S(\mreg/_03865_ ), .Z(\mreg/_01023_ ) );
MUX2_X1 \mreg/_10762_ ( .A(\mreg/_04668_ ), .B(\mreg/_04961_ ), .S(\mreg/_03865_ ), .Z(\mreg/_01024_ ) );
MUX2_X1 \mreg/_10763_ ( .A(\mreg/_04671_ ), .B(\mreg/_04964_ ), .S(\mreg/_03865_ ), .Z(\mreg/_01025_ ) );
MUX2_X1 \mreg/_10764_ ( .A(\mreg/_04672_ ), .B(\mreg/_04965_ ), .S(\mreg/_03865_ ), .Z(\mreg/_01026_ ) );
MUX2_X1 \mreg/_10765_ ( .A(\mreg/_04673_ ), .B(\mreg/_04966_ ), .S(\mreg/_03865_ ), .Z(\mreg/_01027_ ) );
MUX2_X1 \mreg/_10766_ ( .A(\mreg/_04674_ ), .B(\mreg/_04967_ ), .S(\mreg/_03865_ ), .Z(\mreg/_01028_ ) );
MUX2_X1 \mreg/_10767_ ( .A(\mreg/_04675_ ), .B(\mreg/_04968_ ), .S(\mreg/_03865_ ), .Z(\mreg/_01029_ ) );
MUX2_X1 \mreg/_10768_ ( .A(\mreg/_04676_ ), .B(\mreg/_04969_ ), .S(\mreg/_03865_ ), .Z(\mreg/_01030_ ) );
MUX2_X1 \mreg/_10769_ ( .A(\mreg/_04677_ ), .B(\mreg/_04970_ ), .S(\mreg/_03865_ ), .Z(\mreg/_01031_ ) );
BUF_X4 \mreg/_10770_ ( .A(\mreg/_03864_ ), .Z(\mreg/_03866_ ) );
MUX2_X1 \mreg/_10771_ ( .A(\mreg/_04647_ ), .B(\mreg/_04940_ ), .S(\mreg/_03866_ ), .Z(\mreg/_01032_ ) );
MUX2_X1 \mreg/_10772_ ( .A(\mreg/_04648_ ), .B(\mreg/_04941_ ), .S(\mreg/_03866_ ), .Z(\mreg/_01033_ ) );
MUX2_X1 \mreg/_10773_ ( .A(\mreg/_04649_ ), .B(\mreg/_04942_ ), .S(\mreg/_03866_ ), .Z(\mreg/_01034_ ) );
MUX2_X1 \mreg/_10774_ ( .A(\mreg/_04650_ ), .B(\mreg/_04943_ ), .S(\mreg/_03866_ ), .Z(\mreg/_01035_ ) );
MUX2_X1 \mreg/_10775_ ( .A(\mreg/_04651_ ), .B(\mreg/_04944_ ), .S(\mreg/_03866_ ), .Z(\mreg/_01036_ ) );
MUX2_X1 \mreg/_10776_ ( .A(\mreg/_04652_ ), .B(\mreg/_04945_ ), .S(\mreg/_03866_ ), .Z(\mreg/_01037_ ) );
MUX2_X1 \mreg/_10777_ ( .A(\mreg/_04653_ ), .B(\mreg/_04946_ ), .S(\mreg/_03866_ ), .Z(\mreg/_01038_ ) );
MUX2_X1 \mreg/_10778_ ( .A(\mreg/_04654_ ), .B(\mreg/_04947_ ), .S(\mreg/_03866_ ), .Z(\mreg/_01039_ ) );
MUX2_X1 \mreg/_10779_ ( .A(\mreg/_04655_ ), .B(\mreg/_04948_ ), .S(\mreg/_03866_ ), .Z(\mreg/_01040_ ) );
MUX2_X1 \mreg/_10780_ ( .A(\mreg/_04656_ ), .B(\mreg/_04949_ ), .S(\mreg/_03866_ ), .Z(\mreg/_01041_ ) );
BUF_X4 \mreg/_10781_ ( .A(\mreg/_03864_ ), .Z(\mreg/_03867_ ) );
MUX2_X1 \mreg/_10782_ ( .A(\mreg/_04658_ ), .B(\mreg/_04951_ ), .S(\mreg/_03867_ ), .Z(\mreg/_01042_ ) );
MUX2_X1 \mreg/_10783_ ( .A(\mreg/_04659_ ), .B(\mreg/_04952_ ), .S(\mreg/_03867_ ), .Z(\mreg/_01043_ ) );
MUX2_X1 \mreg/_10784_ ( .A(\mreg/_04660_ ), .B(\mreg/_04953_ ), .S(\mreg/_03867_ ), .Z(\mreg/_01044_ ) );
MUX2_X1 \mreg/_10785_ ( .A(\mreg/_04661_ ), .B(\mreg/_04954_ ), .S(\mreg/_03867_ ), .Z(\mreg/_01045_ ) );
MUX2_X1 \mreg/_10786_ ( .A(\mreg/_04662_ ), .B(\mreg/_04955_ ), .S(\mreg/_03867_ ), .Z(\mreg/_01046_ ) );
MUX2_X1 \mreg/_10787_ ( .A(\mreg/_04663_ ), .B(\mreg/_04956_ ), .S(\mreg/_03867_ ), .Z(\mreg/_01047_ ) );
MUX2_X1 \mreg/_10788_ ( .A(\mreg/_04664_ ), .B(\mreg/_04957_ ), .S(\mreg/_03867_ ), .Z(\mreg/_01048_ ) );
MUX2_X1 \mreg/_10789_ ( .A(\mreg/_04665_ ), .B(\mreg/_04958_ ), .S(\mreg/_03867_ ), .Z(\mreg/_01049_ ) );
MUX2_X1 \mreg/_10790_ ( .A(\mreg/_04666_ ), .B(\mreg/_04959_ ), .S(\mreg/_03867_ ), .Z(\mreg/_01050_ ) );
MUX2_X1 \mreg/_10791_ ( .A(\mreg/_04667_ ), .B(\mreg/_04960_ ), .S(\mreg/_03867_ ), .Z(\mreg/_01051_ ) );
MUX2_X1 \mreg/_10792_ ( .A(\mreg/_04669_ ), .B(\mreg/_04962_ ), .S(\mreg/_03864_ ), .Z(\mreg/_01052_ ) );
MUX2_X1 \mreg/_10793_ ( .A(\mreg/_04670_ ), .B(\mreg/_04963_ ), .S(\mreg/_03864_ ), .Z(\mreg/_01053_ ) );
DFF_X1 \mreg/_10794_ ( .CK(clk ), .D(\mreg/_05933_ ), .Q(\mreg/rf[31][0] ), .QN(\mreg/_05932_ ) );
DFF_X1 \mreg/_10795_ ( .CK(clk ), .D(\mreg/_05934_ ), .Q(\mreg/rf[31][1] ), .QN(\mreg/_00000_ ) );
DFF_X1 \mreg/_10796_ ( .CK(clk ), .D(\mreg/_05935_ ), .Q(\mreg/rf[31][2] ), .QN(\mreg/_00001_ ) );
DFF_X1 \mreg/_10797_ ( .CK(clk ), .D(\mreg/_05936_ ), .Q(\mreg/rf[31][3] ), .QN(\mreg/_00002_ ) );
DFF_X1 \mreg/_10798_ ( .CK(clk ), .D(\mreg/_05937_ ), .Q(\mreg/rf[31][4] ), .QN(\mreg/_00003_ ) );
DFF_X1 \mreg/_10799_ ( .CK(clk ), .D(\mreg/_05938_ ), .Q(\mreg/rf[31][5] ), .QN(\mreg/_00004_ ) );
DFF_X1 \mreg/_10800_ ( .CK(clk ), .D(\mreg/_05939_ ), .Q(\mreg/rf[31][6] ), .QN(\mreg/_00005_ ) );
DFF_X1 \mreg/_10801_ ( .CK(clk ), .D(\mreg/_05940_ ), .Q(\mreg/rf[31][7] ), .QN(\mreg/_00006_ ) );
DFF_X1 \mreg/_10802_ ( .CK(clk ), .D(\mreg/_05941_ ), .Q(\mreg/rf[31][8] ), .QN(\mreg/_00007_ ) );
DFF_X1 \mreg/_10803_ ( .CK(clk ), .D(\mreg/_05942_ ), .Q(\mreg/rf[31][9] ), .QN(\mreg/_00008_ ) );
DFF_X1 \mreg/_10804_ ( .CK(clk ), .D(\mreg/_05943_ ), .Q(\mreg/rf[31][10] ), .QN(\mreg/_00009_ ) );
DFF_X1 \mreg/_10805_ ( .CK(clk ), .D(\mreg/_05944_ ), .Q(\mreg/rf[31][11] ), .QN(\mreg/_00010_ ) );
DFF_X1 \mreg/_10806_ ( .CK(clk ), .D(\mreg/_05945_ ), .Q(\mreg/rf[31][12] ), .QN(\mreg/_00011_ ) );
DFF_X1 \mreg/_10807_ ( .CK(clk ), .D(\mreg/_05946_ ), .Q(\mreg/rf[31][13] ), .QN(\mreg/_00012_ ) );
DFF_X1 \mreg/_10808_ ( .CK(clk ), .D(\mreg/_05947_ ), .Q(\mreg/rf[31][14] ), .QN(\mreg/_00013_ ) );
DFF_X1 \mreg/_10809_ ( .CK(clk ), .D(\mreg/_05948_ ), .Q(\mreg/rf[31][15] ), .QN(\mreg/_00014_ ) );
DFF_X1 \mreg/_10810_ ( .CK(clk ), .D(\mreg/_05949_ ), .Q(\mreg/rf[31][16] ), .QN(\mreg/_00015_ ) );
DFF_X1 \mreg/_10811_ ( .CK(clk ), .D(\mreg/_05950_ ), .Q(\mreg/rf[31][17] ), .QN(\mreg/_00016_ ) );
DFF_X1 \mreg/_10812_ ( .CK(clk ), .D(\mreg/_05951_ ), .Q(\mreg/rf[31][18] ), .QN(\mreg/_00017_ ) );
DFF_X1 \mreg/_10813_ ( .CK(clk ), .D(\mreg/_05952_ ), .Q(\mreg/rf[31][19] ), .QN(\mreg/_00018_ ) );
DFF_X1 \mreg/_10814_ ( .CK(clk ), .D(\mreg/_05953_ ), .Q(\mreg/rf[31][20] ), .QN(\mreg/_00019_ ) );
DFF_X1 \mreg/_10815_ ( .CK(clk ), .D(\mreg/_05954_ ), .Q(\mreg/rf[31][21] ), .QN(\mreg/_00020_ ) );
DFF_X1 \mreg/_10816_ ( .CK(clk ), .D(\mreg/_05955_ ), .Q(\mreg/rf[31][22] ), .QN(\mreg/_00021_ ) );
DFF_X1 \mreg/_10817_ ( .CK(clk ), .D(\mreg/_05956_ ), .Q(\mreg/rf[31][23] ), .QN(\mreg/_00022_ ) );
DFF_X1 \mreg/_10818_ ( .CK(clk ), .D(\mreg/_05957_ ), .Q(\mreg/rf[31][24] ), .QN(\mreg/_00023_ ) );
DFF_X1 \mreg/_10819_ ( .CK(clk ), .D(\mreg/_05958_ ), .Q(\mreg/rf[31][25] ), .QN(\mreg/_00024_ ) );
DFF_X1 \mreg/_10820_ ( .CK(clk ), .D(\mreg/_05959_ ), .Q(\mreg/rf[31][26] ), .QN(\mreg/_00025_ ) );
DFF_X1 \mreg/_10821_ ( .CK(clk ), .D(\mreg/_05960_ ), .Q(\mreg/rf[31][27] ), .QN(\mreg/_00026_ ) );
DFF_X1 \mreg/_10822_ ( .CK(clk ), .D(\mreg/_05961_ ), .Q(\mreg/rf[31][28] ), .QN(\mreg/_00027_ ) );
DFF_X1 \mreg/_10823_ ( .CK(clk ), .D(\mreg/_05962_ ), .Q(\mreg/rf[31][29] ), .QN(\mreg/_00028_ ) );
DFF_X1 \mreg/_10824_ ( .CK(clk ), .D(\mreg/_05963_ ), .Q(\mreg/rf[31][30] ), .QN(\mreg/_00029_ ) );
DFF_X1 \mreg/_10825_ ( .CK(clk ), .D(\mreg/_05964_ ), .Q(\mreg/rf[31][31] ), .QN(\mreg/_00030_ ) );
DFF_X1 \mreg/_10826_ ( .CK(clk ), .D(\mreg/_05965_ ), .Q(\mreg/rf[1][0] ), .QN(\mreg/_05931_ ) );
DFF_X1 \mreg/_10827_ ( .CK(clk ), .D(\mreg/_05966_ ), .Q(\mreg/rf[1][1] ), .QN(\mreg/_05930_ ) );
DFF_X1 \mreg/_10828_ ( .CK(clk ), .D(\mreg/_05967_ ), .Q(\mreg/rf[1][2] ), .QN(\mreg/_05929_ ) );
DFF_X1 \mreg/_10829_ ( .CK(clk ), .D(\mreg/_05968_ ), .Q(\mreg/rf[1][3] ), .QN(\mreg/_05928_ ) );
DFF_X1 \mreg/_10830_ ( .CK(clk ), .D(\mreg/_05969_ ), .Q(\mreg/rf[1][4] ), .QN(\mreg/_05927_ ) );
DFF_X1 \mreg/_10831_ ( .CK(clk ), .D(\mreg/_05970_ ), .Q(\mreg/rf[1][5] ), .QN(\mreg/_05926_ ) );
DFF_X1 \mreg/_10832_ ( .CK(clk ), .D(\mreg/_05971_ ), .Q(\mreg/rf[1][6] ), .QN(\mreg/_05925_ ) );
DFF_X1 \mreg/_10833_ ( .CK(clk ), .D(\mreg/_05972_ ), .Q(\mreg/rf[1][7] ), .QN(\mreg/_05924_ ) );
DFF_X1 \mreg/_10834_ ( .CK(clk ), .D(\mreg/_05973_ ), .Q(\mreg/rf[1][8] ), .QN(\mreg/_05923_ ) );
DFF_X1 \mreg/_10835_ ( .CK(clk ), .D(\mreg/_05974_ ), .Q(\mreg/rf[1][9] ), .QN(\mreg/_05922_ ) );
DFF_X1 \mreg/_10836_ ( .CK(clk ), .D(\mreg/_05975_ ), .Q(\mreg/rf[1][10] ), .QN(\mreg/_05921_ ) );
DFF_X1 \mreg/_10837_ ( .CK(clk ), .D(\mreg/_05976_ ), .Q(\mreg/rf[1][11] ), .QN(\mreg/_05920_ ) );
DFF_X1 \mreg/_10838_ ( .CK(clk ), .D(\mreg/_05977_ ), .Q(\mreg/rf[1][12] ), .QN(\mreg/_05919_ ) );
DFF_X1 \mreg/_10839_ ( .CK(clk ), .D(\mreg/_05978_ ), .Q(\mreg/rf[1][13] ), .QN(\mreg/_05918_ ) );
DFF_X1 \mreg/_10840_ ( .CK(clk ), .D(\mreg/_05979_ ), .Q(\mreg/rf[1][14] ), .QN(\mreg/_05917_ ) );
DFF_X1 \mreg/_10841_ ( .CK(clk ), .D(\mreg/_05980_ ), .Q(\mreg/rf[1][15] ), .QN(\mreg/_05916_ ) );
DFF_X1 \mreg/_10842_ ( .CK(clk ), .D(\mreg/_05981_ ), .Q(\mreg/rf[1][16] ), .QN(\mreg/_05915_ ) );
DFF_X1 \mreg/_10843_ ( .CK(clk ), .D(\mreg/_05982_ ), .Q(\mreg/rf[1][17] ), .QN(\mreg/_05914_ ) );
DFF_X1 \mreg/_10844_ ( .CK(clk ), .D(\mreg/_05983_ ), .Q(\mreg/rf[1][18] ), .QN(\mreg/_05913_ ) );
DFF_X1 \mreg/_10845_ ( .CK(clk ), .D(\mreg/_05984_ ), .Q(\mreg/rf[1][19] ), .QN(\mreg/_05912_ ) );
DFF_X1 \mreg/_10846_ ( .CK(clk ), .D(\mreg/_05985_ ), .Q(\mreg/rf[1][20] ), .QN(\mreg/_05911_ ) );
DFF_X1 \mreg/_10847_ ( .CK(clk ), .D(\mreg/_05986_ ), .Q(\mreg/rf[1][21] ), .QN(\mreg/_05910_ ) );
DFF_X1 \mreg/_10848_ ( .CK(clk ), .D(\mreg/_05987_ ), .Q(\mreg/rf[1][22] ), .QN(\mreg/_05909_ ) );
DFF_X1 \mreg/_10849_ ( .CK(clk ), .D(\mreg/_05988_ ), .Q(\mreg/rf[1][23] ), .QN(\mreg/_05908_ ) );
DFF_X1 \mreg/_10850_ ( .CK(clk ), .D(\mreg/_05989_ ), .Q(\mreg/rf[1][24] ), .QN(\mreg/_05907_ ) );
DFF_X1 \mreg/_10851_ ( .CK(clk ), .D(\mreg/_05990_ ), .Q(\mreg/rf[1][25] ), .QN(\mreg/_05906_ ) );
DFF_X1 \mreg/_10852_ ( .CK(clk ), .D(\mreg/_05991_ ), .Q(\mreg/rf[1][26] ), .QN(\mreg/_05905_ ) );
DFF_X1 \mreg/_10853_ ( .CK(clk ), .D(\mreg/_05992_ ), .Q(\mreg/rf[1][27] ), .QN(\mreg/_05904_ ) );
DFF_X1 \mreg/_10854_ ( .CK(clk ), .D(\mreg/_05993_ ), .Q(\mreg/rf[1][28] ), .QN(\mreg/_05903_ ) );
DFF_X1 \mreg/_10855_ ( .CK(clk ), .D(\mreg/_05994_ ), .Q(\mreg/rf[1][29] ), .QN(\mreg/_05902_ ) );
DFF_X1 \mreg/_10856_ ( .CK(clk ), .D(\mreg/_05995_ ), .Q(\mreg/rf[1][30] ), .QN(\mreg/_05901_ ) );
DFF_X1 \mreg/_10857_ ( .CK(clk ), .D(\mreg/_05996_ ), .Q(\mreg/rf[1][31] ), .QN(\mreg/_05900_ ) );
DFF_X1 \mreg/_10858_ ( .CK(clk ), .D(\mreg/_05997_ ), .Q(\mreg/rf[2][0] ), .QN(\mreg/_05899_ ) );
DFF_X1 \mreg/_10859_ ( .CK(clk ), .D(\mreg/_05998_ ), .Q(\mreg/rf[2][1] ), .QN(\mreg/_05898_ ) );
DFF_X1 \mreg/_10860_ ( .CK(clk ), .D(\mreg/_05999_ ), .Q(\mreg/rf[2][2] ), .QN(\mreg/_05897_ ) );
DFF_X1 \mreg/_10861_ ( .CK(clk ), .D(\mreg/_06000_ ), .Q(\mreg/rf[2][3] ), .QN(\mreg/_05896_ ) );
DFF_X1 \mreg/_10862_ ( .CK(clk ), .D(\mreg/_06001_ ), .Q(\mreg/rf[2][4] ), .QN(\mreg/_05895_ ) );
DFF_X1 \mreg/_10863_ ( .CK(clk ), .D(\mreg/_06002_ ), .Q(\mreg/rf[2][5] ), .QN(\mreg/_05894_ ) );
DFF_X1 \mreg/_10864_ ( .CK(clk ), .D(\mreg/_06003_ ), .Q(\mreg/rf[2][6] ), .QN(\mreg/_05893_ ) );
DFF_X1 \mreg/_10865_ ( .CK(clk ), .D(\mreg/_06004_ ), .Q(\mreg/rf[2][7] ), .QN(\mreg/_05892_ ) );
DFF_X1 \mreg/_10866_ ( .CK(clk ), .D(\mreg/_06005_ ), .Q(\mreg/rf[2][8] ), .QN(\mreg/_05891_ ) );
DFF_X1 \mreg/_10867_ ( .CK(clk ), .D(\mreg/_06006_ ), .Q(\mreg/rf[2][9] ), .QN(\mreg/_05890_ ) );
DFF_X1 \mreg/_10868_ ( .CK(clk ), .D(\mreg/_06007_ ), .Q(\mreg/rf[2][10] ), .QN(\mreg/_05889_ ) );
DFF_X1 \mreg/_10869_ ( .CK(clk ), .D(\mreg/_06008_ ), .Q(\mreg/rf[2][11] ), .QN(\mreg/_05888_ ) );
DFF_X1 \mreg/_10870_ ( .CK(clk ), .D(\mreg/_06009_ ), .Q(\mreg/rf[2][12] ), .QN(\mreg/_05887_ ) );
DFF_X1 \mreg/_10871_ ( .CK(clk ), .D(\mreg/_06010_ ), .Q(\mreg/rf[2][13] ), .QN(\mreg/_05886_ ) );
DFF_X1 \mreg/_10872_ ( .CK(clk ), .D(\mreg/_06011_ ), .Q(\mreg/rf[2][14] ), .QN(\mreg/_05885_ ) );
DFF_X1 \mreg/_10873_ ( .CK(clk ), .D(\mreg/_06012_ ), .Q(\mreg/rf[2][15] ), .QN(\mreg/_05884_ ) );
DFF_X1 \mreg/_10874_ ( .CK(clk ), .D(\mreg/_06013_ ), .Q(\mreg/rf[2][16] ), .QN(\mreg/_05883_ ) );
DFF_X1 \mreg/_10875_ ( .CK(clk ), .D(\mreg/_06014_ ), .Q(\mreg/rf[2][17] ), .QN(\mreg/_05882_ ) );
DFF_X1 \mreg/_10876_ ( .CK(clk ), .D(\mreg/_06015_ ), .Q(\mreg/rf[2][18] ), .QN(\mreg/_05881_ ) );
DFF_X1 \mreg/_10877_ ( .CK(clk ), .D(\mreg/_06016_ ), .Q(\mreg/rf[2][19] ), .QN(\mreg/_05880_ ) );
DFF_X1 \mreg/_10878_ ( .CK(clk ), .D(\mreg/_06017_ ), .Q(\mreg/rf[2][20] ), .QN(\mreg/_05879_ ) );
DFF_X1 \mreg/_10879_ ( .CK(clk ), .D(\mreg/_06018_ ), .Q(\mreg/rf[2][21] ), .QN(\mreg/_05878_ ) );
DFF_X1 \mreg/_10880_ ( .CK(clk ), .D(\mreg/_06019_ ), .Q(\mreg/rf[2][22] ), .QN(\mreg/_05877_ ) );
DFF_X1 \mreg/_10881_ ( .CK(clk ), .D(\mreg/_06020_ ), .Q(\mreg/rf[2][23] ), .QN(\mreg/_05876_ ) );
DFF_X1 \mreg/_10882_ ( .CK(clk ), .D(\mreg/_06021_ ), .Q(\mreg/rf[2][24] ), .QN(\mreg/_05875_ ) );
DFF_X1 \mreg/_10883_ ( .CK(clk ), .D(\mreg/_06022_ ), .Q(\mreg/rf[2][25] ), .QN(\mreg/_05874_ ) );
DFF_X1 \mreg/_10884_ ( .CK(clk ), .D(\mreg/_06023_ ), .Q(\mreg/rf[2][26] ), .QN(\mreg/_05873_ ) );
DFF_X1 \mreg/_10885_ ( .CK(clk ), .D(\mreg/_06024_ ), .Q(\mreg/rf[2][27] ), .QN(\mreg/_05872_ ) );
DFF_X1 \mreg/_10886_ ( .CK(clk ), .D(\mreg/_06025_ ), .Q(\mreg/rf[2][28] ), .QN(\mreg/_05871_ ) );
DFF_X1 \mreg/_10887_ ( .CK(clk ), .D(\mreg/_06026_ ), .Q(\mreg/rf[2][29] ), .QN(\mreg/_05870_ ) );
DFF_X1 \mreg/_10888_ ( .CK(clk ), .D(\mreg/_06027_ ), .Q(\mreg/rf[2][30] ), .QN(\mreg/_05869_ ) );
DFF_X1 \mreg/_10889_ ( .CK(clk ), .D(\mreg/_06028_ ), .Q(\mreg/rf[2][31] ), .QN(\mreg/_05868_ ) );
DFF_X1 \mreg/_10890_ ( .CK(clk ), .D(\mreg/_06029_ ), .Q(\mreg/rf[3][0] ), .QN(\mreg/_05867_ ) );
DFF_X1 \mreg/_10891_ ( .CK(clk ), .D(\mreg/_06030_ ), .Q(\mreg/rf[3][1] ), .QN(\mreg/_05866_ ) );
DFF_X1 \mreg/_10892_ ( .CK(clk ), .D(\mreg/_06031_ ), .Q(\mreg/rf[3][2] ), .QN(\mreg/_05865_ ) );
DFF_X1 \mreg/_10893_ ( .CK(clk ), .D(\mreg/_06032_ ), .Q(\mreg/rf[3][3] ), .QN(\mreg/_05864_ ) );
DFF_X1 \mreg/_10894_ ( .CK(clk ), .D(\mreg/_06033_ ), .Q(\mreg/rf[3][4] ), .QN(\mreg/_05863_ ) );
DFF_X1 \mreg/_10895_ ( .CK(clk ), .D(\mreg/_06034_ ), .Q(\mreg/rf[3][5] ), .QN(\mreg/_05862_ ) );
DFF_X1 \mreg/_10896_ ( .CK(clk ), .D(\mreg/_06035_ ), .Q(\mreg/rf[3][6] ), .QN(\mreg/_05861_ ) );
DFF_X1 \mreg/_10897_ ( .CK(clk ), .D(\mreg/_06036_ ), .Q(\mreg/rf[3][7] ), .QN(\mreg/_05860_ ) );
DFF_X1 \mreg/_10898_ ( .CK(clk ), .D(\mreg/_06037_ ), .Q(\mreg/rf[3][8] ), .QN(\mreg/_05859_ ) );
DFF_X1 \mreg/_10899_ ( .CK(clk ), .D(\mreg/_06038_ ), .Q(\mreg/rf[3][9] ), .QN(\mreg/_05858_ ) );
DFF_X1 \mreg/_10900_ ( .CK(clk ), .D(\mreg/_06039_ ), .Q(\mreg/rf[3][10] ), .QN(\mreg/_05857_ ) );
DFF_X1 \mreg/_10901_ ( .CK(clk ), .D(\mreg/_06040_ ), .Q(\mreg/rf[3][11] ), .QN(\mreg/_05856_ ) );
DFF_X1 \mreg/_10902_ ( .CK(clk ), .D(\mreg/_06041_ ), .Q(\mreg/rf[3][12] ), .QN(\mreg/_05855_ ) );
DFF_X1 \mreg/_10903_ ( .CK(clk ), .D(\mreg/_06042_ ), .Q(\mreg/rf[3][13] ), .QN(\mreg/_05854_ ) );
DFF_X1 \mreg/_10904_ ( .CK(clk ), .D(\mreg/_06043_ ), .Q(\mreg/rf[3][14] ), .QN(\mreg/_05853_ ) );
DFF_X1 \mreg/_10905_ ( .CK(clk ), .D(\mreg/_06044_ ), .Q(\mreg/rf[3][15] ), .QN(\mreg/_05852_ ) );
DFF_X1 \mreg/_10906_ ( .CK(clk ), .D(\mreg/_06045_ ), .Q(\mreg/rf[3][16] ), .QN(\mreg/_05851_ ) );
DFF_X1 \mreg/_10907_ ( .CK(clk ), .D(\mreg/_06046_ ), .Q(\mreg/rf[3][17] ), .QN(\mreg/_05850_ ) );
DFF_X1 \mreg/_10908_ ( .CK(clk ), .D(\mreg/_06047_ ), .Q(\mreg/rf[3][18] ), .QN(\mreg/_05849_ ) );
DFF_X1 \mreg/_10909_ ( .CK(clk ), .D(\mreg/_06048_ ), .Q(\mreg/rf[3][19] ), .QN(\mreg/_05848_ ) );
DFF_X1 \mreg/_10910_ ( .CK(clk ), .D(\mreg/_06049_ ), .Q(\mreg/rf[3][20] ), .QN(\mreg/_05847_ ) );
DFF_X1 \mreg/_10911_ ( .CK(clk ), .D(\mreg/_06050_ ), .Q(\mreg/rf[3][21] ), .QN(\mreg/_05846_ ) );
DFF_X1 \mreg/_10912_ ( .CK(clk ), .D(\mreg/_06051_ ), .Q(\mreg/rf[3][22] ), .QN(\mreg/_05845_ ) );
DFF_X1 \mreg/_10913_ ( .CK(clk ), .D(\mreg/_06052_ ), .Q(\mreg/rf[3][23] ), .QN(\mreg/_05844_ ) );
DFF_X1 \mreg/_10914_ ( .CK(clk ), .D(\mreg/_06053_ ), .Q(\mreg/rf[3][24] ), .QN(\mreg/_05843_ ) );
DFF_X1 \mreg/_10915_ ( .CK(clk ), .D(\mreg/_06054_ ), .Q(\mreg/rf[3][25] ), .QN(\mreg/_05842_ ) );
DFF_X1 \mreg/_10916_ ( .CK(clk ), .D(\mreg/_06055_ ), .Q(\mreg/rf[3][26] ), .QN(\mreg/_05841_ ) );
DFF_X1 \mreg/_10917_ ( .CK(clk ), .D(\mreg/_06056_ ), .Q(\mreg/rf[3][27] ), .QN(\mreg/_05840_ ) );
DFF_X1 \mreg/_10918_ ( .CK(clk ), .D(\mreg/_06057_ ), .Q(\mreg/rf[3][28] ), .QN(\mreg/_05839_ ) );
DFF_X1 \mreg/_10919_ ( .CK(clk ), .D(\mreg/_06058_ ), .Q(\mreg/rf[3][29] ), .QN(\mreg/_05838_ ) );
DFF_X1 \mreg/_10920_ ( .CK(clk ), .D(\mreg/_06059_ ), .Q(\mreg/rf[3][30] ), .QN(\mreg/_05837_ ) );
DFF_X1 \mreg/_10921_ ( .CK(clk ), .D(\mreg/_06060_ ), .Q(\mreg/rf[3][31] ), .QN(\mreg/_05836_ ) );
DFF_X1 \mreg/_10922_ ( .CK(clk ), .D(\mreg/_06061_ ), .Q(\mreg/rf[4][0] ), .QN(\mreg/_05835_ ) );
DFF_X1 \mreg/_10923_ ( .CK(clk ), .D(\mreg/_06062_ ), .Q(\mreg/rf[4][1] ), .QN(\mreg/_05834_ ) );
DFF_X1 \mreg/_10924_ ( .CK(clk ), .D(\mreg/_06063_ ), .Q(\mreg/rf[4][2] ), .QN(\mreg/_05833_ ) );
DFF_X1 \mreg/_10925_ ( .CK(clk ), .D(\mreg/_06064_ ), .Q(\mreg/rf[4][3] ), .QN(\mreg/_05832_ ) );
DFF_X1 \mreg/_10926_ ( .CK(clk ), .D(\mreg/_06065_ ), .Q(\mreg/rf[4][4] ), .QN(\mreg/_05831_ ) );
DFF_X1 \mreg/_10927_ ( .CK(clk ), .D(\mreg/_06066_ ), .Q(\mreg/rf[4][5] ), .QN(\mreg/_05830_ ) );
DFF_X1 \mreg/_10928_ ( .CK(clk ), .D(\mreg/_06067_ ), .Q(\mreg/rf[4][6] ), .QN(\mreg/_05829_ ) );
DFF_X1 \mreg/_10929_ ( .CK(clk ), .D(\mreg/_06068_ ), .Q(\mreg/rf[4][7] ), .QN(\mreg/_05828_ ) );
DFF_X1 \mreg/_10930_ ( .CK(clk ), .D(\mreg/_06069_ ), .Q(\mreg/rf[4][8] ), .QN(\mreg/_05827_ ) );
DFF_X1 \mreg/_10931_ ( .CK(clk ), .D(\mreg/_06070_ ), .Q(\mreg/rf[4][9] ), .QN(\mreg/_05826_ ) );
DFF_X1 \mreg/_10932_ ( .CK(clk ), .D(\mreg/_06071_ ), .Q(\mreg/rf[4][10] ), .QN(\mreg/_05825_ ) );
DFF_X1 \mreg/_10933_ ( .CK(clk ), .D(\mreg/_06072_ ), .Q(\mreg/rf[4][11] ), .QN(\mreg/_05824_ ) );
DFF_X1 \mreg/_10934_ ( .CK(clk ), .D(\mreg/_06073_ ), .Q(\mreg/rf[4][12] ), .QN(\mreg/_05823_ ) );
DFF_X1 \mreg/_10935_ ( .CK(clk ), .D(\mreg/_06074_ ), .Q(\mreg/rf[4][13] ), .QN(\mreg/_05822_ ) );
DFF_X1 \mreg/_10936_ ( .CK(clk ), .D(\mreg/_06075_ ), .Q(\mreg/rf[4][14] ), .QN(\mreg/_05821_ ) );
DFF_X1 \mreg/_10937_ ( .CK(clk ), .D(\mreg/_06076_ ), .Q(\mreg/rf[4][15] ), .QN(\mreg/_05820_ ) );
DFF_X1 \mreg/_10938_ ( .CK(clk ), .D(\mreg/_06077_ ), .Q(\mreg/rf[4][16] ), .QN(\mreg/_05819_ ) );
DFF_X1 \mreg/_10939_ ( .CK(clk ), .D(\mreg/_06078_ ), .Q(\mreg/rf[4][17] ), .QN(\mreg/_05818_ ) );
DFF_X1 \mreg/_10940_ ( .CK(clk ), .D(\mreg/_06079_ ), .Q(\mreg/rf[4][18] ), .QN(\mreg/_05817_ ) );
DFF_X1 \mreg/_10941_ ( .CK(clk ), .D(\mreg/_06080_ ), .Q(\mreg/rf[4][19] ), .QN(\mreg/_05816_ ) );
DFF_X1 \mreg/_10942_ ( .CK(clk ), .D(\mreg/_06081_ ), .Q(\mreg/rf[4][20] ), .QN(\mreg/_05815_ ) );
DFF_X1 \mreg/_10943_ ( .CK(clk ), .D(\mreg/_06082_ ), .Q(\mreg/rf[4][21] ), .QN(\mreg/_05814_ ) );
DFF_X1 \mreg/_10944_ ( .CK(clk ), .D(\mreg/_06083_ ), .Q(\mreg/rf[4][22] ), .QN(\mreg/_05813_ ) );
DFF_X1 \mreg/_10945_ ( .CK(clk ), .D(\mreg/_06084_ ), .Q(\mreg/rf[4][23] ), .QN(\mreg/_05812_ ) );
DFF_X1 \mreg/_10946_ ( .CK(clk ), .D(\mreg/_06085_ ), .Q(\mreg/rf[4][24] ), .QN(\mreg/_05811_ ) );
DFF_X1 \mreg/_10947_ ( .CK(clk ), .D(\mreg/_06086_ ), .Q(\mreg/rf[4][25] ), .QN(\mreg/_05810_ ) );
DFF_X1 \mreg/_10948_ ( .CK(clk ), .D(\mreg/_06087_ ), .Q(\mreg/rf[4][26] ), .QN(\mreg/_05809_ ) );
DFF_X1 \mreg/_10949_ ( .CK(clk ), .D(\mreg/_06088_ ), .Q(\mreg/rf[4][27] ), .QN(\mreg/_05808_ ) );
DFF_X1 \mreg/_10950_ ( .CK(clk ), .D(\mreg/_06089_ ), .Q(\mreg/rf[4][28] ), .QN(\mreg/_05807_ ) );
DFF_X1 \mreg/_10951_ ( .CK(clk ), .D(\mreg/_06090_ ), .Q(\mreg/rf[4][29] ), .QN(\mreg/_05806_ ) );
DFF_X1 \mreg/_10952_ ( .CK(clk ), .D(\mreg/_06091_ ), .Q(\mreg/rf[4][30] ), .QN(\mreg/_05805_ ) );
DFF_X1 \mreg/_10953_ ( .CK(clk ), .D(\mreg/_06092_ ), .Q(\mreg/rf[4][31] ), .QN(\mreg/_05804_ ) );
DFF_X1 \mreg/_10954_ ( .CK(clk ), .D(\mreg/_06093_ ), .Q(\mreg/rf[5][0] ), .QN(\mreg/_05803_ ) );
DFF_X1 \mreg/_10955_ ( .CK(clk ), .D(\mreg/_06094_ ), .Q(\mreg/rf[5][1] ), .QN(\mreg/_05802_ ) );
DFF_X1 \mreg/_10956_ ( .CK(clk ), .D(\mreg/_06095_ ), .Q(\mreg/rf[5][2] ), .QN(\mreg/_05801_ ) );
DFF_X1 \mreg/_10957_ ( .CK(clk ), .D(\mreg/_06096_ ), .Q(\mreg/rf[5][3] ), .QN(\mreg/_05800_ ) );
DFF_X1 \mreg/_10958_ ( .CK(clk ), .D(\mreg/_06097_ ), .Q(\mreg/rf[5][4] ), .QN(\mreg/_05799_ ) );
DFF_X1 \mreg/_10959_ ( .CK(clk ), .D(\mreg/_06098_ ), .Q(\mreg/rf[5][5] ), .QN(\mreg/_05798_ ) );
DFF_X1 \mreg/_10960_ ( .CK(clk ), .D(\mreg/_06099_ ), .Q(\mreg/rf[5][6] ), .QN(\mreg/_05797_ ) );
DFF_X1 \mreg/_10961_ ( .CK(clk ), .D(\mreg/_06100_ ), .Q(\mreg/rf[5][7] ), .QN(\mreg/_05796_ ) );
DFF_X1 \mreg/_10962_ ( .CK(clk ), .D(\mreg/_06101_ ), .Q(\mreg/rf[5][8] ), .QN(\mreg/_05795_ ) );
DFF_X1 \mreg/_10963_ ( .CK(clk ), .D(\mreg/_06102_ ), .Q(\mreg/rf[5][9] ), .QN(\mreg/_05794_ ) );
DFF_X1 \mreg/_10964_ ( .CK(clk ), .D(\mreg/_06103_ ), .Q(\mreg/rf[5][10] ), .QN(\mreg/_05793_ ) );
DFF_X1 \mreg/_10965_ ( .CK(clk ), .D(\mreg/_06104_ ), .Q(\mreg/rf[5][11] ), .QN(\mreg/_05792_ ) );
DFF_X1 \mreg/_10966_ ( .CK(clk ), .D(\mreg/_06105_ ), .Q(\mreg/rf[5][12] ), .QN(\mreg/_05791_ ) );
DFF_X1 \mreg/_10967_ ( .CK(clk ), .D(\mreg/_06106_ ), .Q(\mreg/rf[5][13] ), .QN(\mreg/_05790_ ) );
DFF_X1 \mreg/_10968_ ( .CK(clk ), .D(\mreg/_06107_ ), .Q(\mreg/rf[5][14] ), .QN(\mreg/_05789_ ) );
DFF_X1 \mreg/_10969_ ( .CK(clk ), .D(\mreg/_06108_ ), .Q(\mreg/rf[5][15] ), .QN(\mreg/_05788_ ) );
DFF_X1 \mreg/_10970_ ( .CK(clk ), .D(\mreg/_06109_ ), .Q(\mreg/rf[5][16] ), .QN(\mreg/_05787_ ) );
DFF_X1 \mreg/_10971_ ( .CK(clk ), .D(\mreg/_06110_ ), .Q(\mreg/rf[5][17] ), .QN(\mreg/_05786_ ) );
DFF_X1 \mreg/_10972_ ( .CK(clk ), .D(\mreg/_06111_ ), .Q(\mreg/rf[5][18] ), .QN(\mreg/_05785_ ) );
DFF_X1 \mreg/_10973_ ( .CK(clk ), .D(\mreg/_06112_ ), .Q(\mreg/rf[5][19] ), .QN(\mreg/_05784_ ) );
DFF_X1 \mreg/_10974_ ( .CK(clk ), .D(\mreg/_06113_ ), .Q(\mreg/rf[5][20] ), .QN(\mreg/_05783_ ) );
DFF_X1 \mreg/_10975_ ( .CK(clk ), .D(\mreg/_06114_ ), .Q(\mreg/rf[5][21] ), .QN(\mreg/_05782_ ) );
DFF_X1 \mreg/_10976_ ( .CK(clk ), .D(\mreg/_06115_ ), .Q(\mreg/rf[5][22] ), .QN(\mreg/_05781_ ) );
DFF_X1 \mreg/_10977_ ( .CK(clk ), .D(\mreg/_06116_ ), .Q(\mreg/rf[5][23] ), .QN(\mreg/_05780_ ) );
DFF_X1 \mreg/_10978_ ( .CK(clk ), .D(\mreg/_06117_ ), .Q(\mreg/rf[5][24] ), .QN(\mreg/_05779_ ) );
DFF_X1 \mreg/_10979_ ( .CK(clk ), .D(\mreg/_06118_ ), .Q(\mreg/rf[5][25] ), .QN(\mreg/_05778_ ) );
DFF_X1 \mreg/_10980_ ( .CK(clk ), .D(\mreg/_06119_ ), .Q(\mreg/rf[5][26] ), .QN(\mreg/_05777_ ) );
DFF_X1 \mreg/_10981_ ( .CK(clk ), .D(\mreg/_06120_ ), .Q(\mreg/rf[5][27] ), .QN(\mreg/_05776_ ) );
DFF_X1 \mreg/_10982_ ( .CK(clk ), .D(\mreg/_06121_ ), .Q(\mreg/rf[5][28] ), .QN(\mreg/_05775_ ) );
DFF_X1 \mreg/_10983_ ( .CK(clk ), .D(\mreg/_06122_ ), .Q(\mreg/rf[5][29] ), .QN(\mreg/_05774_ ) );
DFF_X1 \mreg/_10984_ ( .CK(clk ), .D(\mreg/_06123_ ), .Q(\mreg/rf[5][30] ), .QN(\mreg/_05773_ ) );
DFF_X1 \mreg/_10985_ ( .CK(clk ), .D(\mreg/_06124_ ), .Q(\mreg/rf[5][31] ), .QN(\mreg/_05772_ ) );
DFF_X1 \mreg/_10986_ ( .CK(clk ), .D(\mreg/_06125_ ), .Q(\mreg/rf[6][0] ), .QN(\mreg/_05771_ ) );
DFF_X1 \mreg/_10987_ ( .CK(clk ), .D(\mreg/_06126_ ), .Q(\mreg/rf[6][1] ), .QN(\mreg/_05770_ ) );
DFF_X1 \mreg/_10988_ ( .CK(clk ), .D(\mreg/_06127_ ), .Q(\mreg/rf[6][2] ), .QN(\mreg/_05769_ ) );
DFF_X1 \mreg/_10989_ ( .CK(clk ), .D(\mreg/_06128_ ), .Q(\mreg/rf[6][3] ), .QN(\mreg/_05768_ ) );
DFF_X1 \mreg/_10990_ ( .CK(clk ), .D(\mreg/_06129_ ), .Q(\mreg/rf[6][4] ), .QN(\mreg/_05767_ ) );
DFF_X1 \mreg/_10991_ ( .CK(clk ), .D(\mreg/_06130_ ), .Q(\mreg/rf[6][5] ), .QN(\mreg/_05766_ ) );
DFF_X1 \mreg/_10992_ ( .CK(clk ), .D(\mreg/_06131_ ), .Q(\mreg/rf[6][6] ), .QN(\mreg/_05765_ ) );
DFF_X1 \mreg/_10993_ ( .CK(clk ), .D(\mreg/_06132_ ), .Q(\mreg/rf[6][7] ), .QN(\mreg/_05764_ ) );
DFF_X1 \mreg/_10994_ ( .CK(clk ), .D(\mreg/_06133_ ), .Q(\mreg/rf[6][8] ), .QN(\mreg/_05763_ ) );
DFF_X1 \mreg/_10995_ ( .CK(clk ), .D(\mreg/_06134_ ), .Q(\mreg/rf[6][9] ), .QN(\mreg/_05762_ ) );
DFF_X1 \mreg/_10996_ ( .CK(clk ), .D(\mreg/_06135_ ), .Q(\mreg/rf[6][10] ), .QN(\mreg/_05761_ ) );
DFF_X1 \mreg/_10997_ ( .CK(clk ), .D(\mreg/_06136_ ), .Q(\mreg/rf[6][11] ), .QN(\mreg/_05760_ ) );
DFF_X1 \mreg/_10998_ ( .CK(clk ), .D(\mreg/_06137_ ), .Q(\mreg/rf[6][12] ), .QN(\mreg/_05759_ ) );
DFF_X1 \mreg/_10999_ ( .CK(clk ), .D(\mreg/_06138_ ), .Q(\mreg/rf[6][13] ), .QN(\mreg/_05758_ ) );
DFF_X1 \mreg/_11000_ ( .CK(clk ), .D(\mreg/_06139_ ), .Q(\mreg/rf[6][14] ), .QN(\mreg/_05757_ ) );
DFF_X1 \mreg/_11001_ ( .CK(clk ), .D(\mreg/_06140_ ), .Q(\mreg/rf[6][15] ), .QN(\mreg/_05756_ ) );
DFF_X1 \mreg/_11002_ ( .CK(clk ), .D(\mreg/_06141_ ), .Q(\mreg/rf[6][16] ), .QN(\mreg/_05755_ ) );
DFF_X1 \mreg/_11003_ ( .CK(clk ), .D(\mreg/_06142_ ), .Q(\mreg/rf[6][17] ), .QN(\mreg/_05754_ ) );
DFF_X1 \mreg/_11004_ ( .CK(clk ), .D(\mreg/_06143_ ), .Q(\mreg/rf[6][18] ), .QN(\mreg/_05753_ ) );
DFF_X1 \mreg/_11005_ ( .CK(clk ), .D(\mreg/_06144_ ), .Q(\mreg/rf[6][19] ), .QN(\mreg/_05752_ ) );
DFF_X1 \mreg/_11006_ ( .CK(clk ), .D(\mreg/_06145_ ), .Q(\mreg/rf[6][20] ), .QN(\mreg/_05751_ ) );
DFF_X1 \mreg/_11007_ ( .CK(clk ), .D(\mreg/_06146_ ), .Q(\mreg/rf[6][21] ), .QN(\mreg/_05750_ ) );
DFF_X1 \mreg/_11008_ ( .CK(clk ), .D(\mreg/_06147_ ), .Q(\mreg/rf[6][22] ), .QN(\mreg/_05749_ ) );
DFF_X1 \mreg/_11009_ ( .CK(clk ), .D(\mreg/_06148_ ), .Q(\mreg/rf[6][23] ), .QN(\mreg/_05748_ ) );
DFF_X1 \mreg/_11010_ ( .CK(clk ), .D(\mreg/_06149_ ), .Q(\mreg/rf[6][24] ), .QN(\mreg/_05747_ ) );
DFF_X1 \mreg/_11011_ ( .CK(clk ), .D(\mreg/_06150_ ), .Q(\mreg/rf[6][25] ), .QN(\mreg/_05746_ ) );
DFF_X1 \mreg/_11012_ ( .CK(clk ), .D(\mreg/_06151_ ), .Q(\mreg/rf[6][26] ), .QN(\mreg/_05745_ ) );
DFF_X1 \mreg/_11013_ ( .CK(clk ), .D(\mreg/_06152_ ), .Q(\mreg/rf[6][27] ), .QN(\mreg/_05744_ ) );
DFF_X1 \mreg/_11014_ ( .CK(clk ), .D(\mreg/_06153_ ), .Q(\mreg/rf[6][28] ), .QN(\mreg/_05743_ ) );
DFF_X1 \mreg/_11015_ ( .CK(clk ), .D(\mreg/_06154_ ), .Q(\mreg/rf[6][29] ), .QN(\mreg/_05742_ ) );
DFF_X1 \mreg/_11016_ ( .CK(clk ), .D(\mreg/_06155_ ), .Q(\mreg/rf[6][30] ), .QN(\mreg/_05741_ ) );
DFF_X1 \mreg/_11017_ ( .CK(clk ), .D(\mreg/_06156_ ), .Q(\mreg/rf[6][31] ), .QN(\mreg/_05740_ ) );
DFF_X1 \mreg/_11018_ ( .CK(clk ), .D(\mreg/_06157_ ), .Q(\mreg/rf[7][0] ), .QN(\mreg/_05739_ ) );
DFF_X1 \mreg/_11019_ ( .CK(clk ), .D(\mreg/_06158_ ), .Q(\mreg/rf[7][1] ), .QN(\mreg/_05738_ ) );
DFF_X1 \mreg/_11020_ ( .CK(clk ), .D(\mreg/_06159_ ), .Q(\mreg/rf[7][2] ), .QN(\mreg/_05737_ ) );
DFF_X1 \mreg/_11021_ ( .CK(clk ), .D(\mreg/_06160_ ), .Q(\mreg/rf[7][3] ), .QN(\mreg/_05736_ ) );
DFF_X1 \mreg/_11022_ ( .CK(clk ), .D(\mreg/_06161_ ), .Q(\mreg/rf[7][4] ), .QN(\mreg/_05735_ ) );
DFF_X1 \mreg/_11023_ ( .CK(clk ), .D(\mreg/_06162_ ), .Q(\mreg/rf[7][5] ), .QN(\mreg/_05734_ ) );
DFF_X1 \mreg/_11024_ ( .CK(clk ), .D(\mreg/_06163_ ), .Q(\mreg/rf[7][6] ), .QN(\mreg/_05733_ ) );
DFF_X1 \mreg/_11025_ ( .CK(clk ), .D(\mreg/_06164_ ), .Q(\mreg/rf[7][7] ), .QN(\mreg/_05732_ ) );
DFF_X1 \mreg/_11026_ ( .CK(clk ), .D(\mreg/_06165_ ), .Q(\mreg/rf[7][8] ), .QN(\mreg/_05731_ ) );
DFF_X1 \mreg/_11027_ ( .CK(clk ), .D(\mreg/_06166_ ), .Q(\mreg/rf[7][9] ), .QN(\mreg/_05730_ ) );
DFF_X1 \mreg/_11028_ ( .CK(clk ), .D(\mreg/_06167_ ), .Q(\mreg/rf[7][10] ), .QN(\mreg/_05729_ ) );
DFF_X1 \mreg/_11029_ ( .CK(clk ), .D(\mreg/_06168_ ), .Q(\mreg/rf[7][11] ), .QN(\mreg/_05728_ ) );
DFF_X1 \mreg/_11030_ ( .CK(clk ), .D(\mreg/_06169_ ), .Q(\mreg/rf[7][12] ), .QN(\mreg/_05727_ ) );
DFF_X1 \mreg/_11031_ ( .CK(clk ), .D(\mreg/_06170_ ), .Q(\mreg/rf[7][13] ), .QN(\mreg/_05726_ ) );
DFF_X1 \mreg/_11032_ ( .CK(clk ), .D(\mreg/_06171_ ), .Q(\mreg/rf[7][14] ), .QN(\mreg/_05725_ ) );
DFF_X1 \mreg/_11033_ ( .CK(clk ), .D(\mreg/_06172_ ), .Q(\mreg/rf[7][15] ), .QN(\mreg/_05724_ ) );
DFF_X1 \mreg/_11034_ ( .CK(clk ), .D(\mreg/_06173_ ), .Q(\mreg/rf[7][16] ), .QN(\mreg/_05723_ ) );
DFF_X1 \mreg/_11035_ ( .CK(clk ), .D(\mreg/_06174_ ), .Q(\mreg/rf[7][17] ), .QN(\mreg/_05722_ ) );
DFF_X1 \mreg/_11036_ ( .CK(clk ), .D(\mreg/_06175_ ), .Q(\mreg/rf[7][18] ), .QN(\mreg/_05721_ ) );
DFF_X1 \mreg/_11037_ ( .CK(clk ), .D(\mreg/_06176_ ), .Q(\mreg/rf[7][19] ), .QN(\mreg/_05720_ ) );
DFF_X1 \mreg/_11038_ ( .CK(clk ), .D(\mreg/_06177_ ), .Q(\mreg/rf[7][20] ), .QN(\mreg/_05719_ ) );
DFF_X1 \mreg/_11039_ ( .CK(clk ), .D(\mreg/_06178_ ), .Q(\mreg/rf[7][21] ), .QN(\mreg/_05718_ ) );
DFF_X1 \mreg/_11040_ ( .CK(clk ), .D(\mreg/_06179_ ), .Q(\mreg/rf[7][22] ), .QN(\mreg/_05717_ ) );
DFF_X1 \mreg/_11041_ ( .CK(clk ), .D(\mreg/_06180_ ), .Q(\mreg/rf[7][23] ), .QN(\mreg/_05716_ ) );
DFF_X1 \mreg/_11042_ ( .CK(clk ), .D(\mreg/_06181_ ), .Q(\mreg/rf[7][24] ), .QN(\mreg/_05715_ ) );
DFF_X1 \mreg/_11043_ ( .CK(clk ), .D(\mreg/_06182_ ), .Q(\mreg/rf[7][25] ), .QN(\mreg/_05714_ ) );
DFF_X1 \mreg/_11044_ ( .CK(clk ), .D(\mreg/_06183_ ), .Q(\mreg/rf[7][26] ), .QN(\mreg/_05713_ ) );
DFF_X1 \mreg/_11045_ ( .CK(clk ), .D(\mreg/_06184_ ), .Q(\mreg/rf[7][27] ), .QN(\mreg/_05712_ ) );
DFF_X1 \mreg/_11046_ ( .CK(clk ), .D(\mreg/_06185_ ), .Q(\mreg/rf[7][28] ), .QN(\mreg/_05711_ ) );
DFF_X1 \mreg/_11047_ ( .CK(clk ), .D(\mreg/_06186_ ), .Q(\mreg/rf[7][29] ), .QN(\mreg/_05710_ ) );
DFF_X1 \mreg/_11048_ ( .CK(clk ), .D(\mreg/_06187_ ), .Q(\mreg/rf[7][30] ), .QN(\mreg/_05709_ ) );
DFF_X1 \mreg/_11049_ ( .CK(clk ), .D(\mreg/_06188_ ), .Q(\mreg/rf[7][31] ), .QN(\mreg/_05708_ ) );
DFF_X1 \mreg/_11050_ ( .CK(clk ), .D(\mreg/_06189_ ), .Q(\mreg/rf[8][0] ), .QN(\mreg/_05707_ ) );
DFF_X1 \mreg/_11051_ ( .CK(clk ), .D(\mreg/_06190_ ), .Q(\mreg/rf[8][1] ), .QN(\mreg/_05706_ ) );
DFF_X1 \mreg/_11052_ ( .CK(clk ), .D(\mreg/_06191_ ), .Q(\mreg/rf[8][2] ), .QN(\mreg/_05705_ ) );
DFF_X1 \mreg/_11053_ ( .CK(clk ), .D(\mreg/_06192_ ), .Q(\mreg/rf[8][3] ), .QN(\mreg/_05704_ ) );
DFF_X1 \mreg/_11054_ ( .CK(clk ), .D(\mreg/_06193_ ), .Q(\mreg/rf[8][4] ), .QN(\mreg/_05703_ ) );
DFF_X1 \mreg/_11055_ ( .CK(clk ), .D(\mreg/_06194_ ), .Q(\mreg/rf[8][5] ), .QN(\mreg/_05702_ ) );
DFF_X1 \mreg/_11056_ ( .CK(clk ), .D(\mreg/_06195_ ), .Q(\mreg/rf[8][6] ), .QN(\mreg/_05701_ ) );
DFF_X1 \mreg/_11057_ ( .CK(clk ), .D(\mreg/_06196_ ), .Q(\mreg/rf[8][7] ), .QN(\mreg/_05700_ ) );
DFF_X1 \mreg/_11058_ ( .CK(clk ), .D(\mreg/_06197_ ), .Q(\mreg/rf[8][8] ), .QN(\mreg/_05699_ ) );
DFF_X1 \mreg/_11059_ ( .CK(clk ), .D(\mreg/_06198_ ), .Q(\mreg/rf[8][9] ), .QN(\mreg/_05698_ ) );
DFF_X1 \mreg/_11060_ ( .CK(clk ), .D(\mreg/_06199_ ), .Q(\mreg/rf[8][10] ), .QN(\mreg/_05697_ ) );
DFF_X1 \mreg/_11061_ ( .CK(clk ), .D(\mreg/_06200_ ), .Q(\mreg/rf[8][11] ), .QN(\mreg/_05696_ ) );
DFF_X1 \mreg/_11062_ ( .CK(clk ), .D(\mreg/_06201_ ), .Q(\mreg/rf[8][12] ), .QN(\mreg/_05695_ ) );
DFF_X1 \mreg/_11063_ ( .CK(clk ), .D(\mreg/_06202_ ), .Q(\mreg/rf[8][13] ), .QN(\mreg/_05694_ ) );
DFF_X1 \mreg/_11064_ ( .CK(clk ), .D(\mreg/_06203_ ), .Q(\mreg/rf[8][14] ), .QN(\mreg/_05693_ ) );
DFF_X1 \mreg/_11065_ ( .CK(clk ), .D(\mreg/_06204_ ), .Q(\mreg/rf[8][15] ), .QN(\mreg/_05692_ ) );
DFF_X1 \mreg/_11066_ ( .CK(clk ), .D(\mreg/_06205_ ), .Q(\mreg/rf[8][16] ), .QN(\mreg/_05691_ ) );
DFF_X1 \mreg/_11067_ ( .CK(clk ), .D(\mreg/_06206_ ), .Q(\mreg/rf[8][17] ), .QN(\mreg/_05690_ ) );
DFF_X1 \mreg/_11068_ ( .CK(clk ), .D(\mreg/_06207_ ), .Q(\mreg/rf[8][18] ), .QN(\mreg/_05689_ ) );
DFF_X1 \mreg/_11069_ ( .CK(clk ), .D(\mreg/_06208_ ), .Q(\mreg/rf[8][19] ), .QN(\mreg/_05688_ ) );
DFF_X1 \mreg/_11070_ ( .CK(clk ), .D(\mreg/_06209_ ), .Q(\mreg/rf[8][20] ), .QN(\mreg/_05687_ ) );
DFF_X1 \mreg/_11071_ ( .CK(clk ), .D(\mreg/_06210_ ), .Q(\mreg/rf[8][21] ), .QN(\mreg/_05686_ ) );
DFF_X1 \mreg/_11072_ ( .CK(clk ), .D(\mreg/_06211_ ), .Q(\mreg/rf[8][22] ), .QN(\mreg/_05685_ ) );
DFF_X1 \mreg/_11073_ ( .CK(clk ), .D(\mreg/_06212_ ), .Q(\mreg/rf[8][23] ), .QN(\mreg/_05684_ ) );
DFF_X1 \mreg/_11074_ ( .CK(clk ), .D(\mreg/_06213_ ), .Q(\mreg/rf[8][24] ), .QN(\mreg/_05683_ ) );
DFF_X1 \mreg/_11075_ ( .CK(clk ), .D(\mreg/_06214_ ), .Q(\mreg/rf[8][25] ), .QN(\mreg/_05682_ ) );
DFF_X1 \mreg/_11076_ ( .CK(clk ), .D(\mreg/_06215_ ), .Q(\mreg/rf[8][26] ), .QN(\mreg/_05681_ ) );
DFF_X1 \mreg/_11077_ ( .CK(clk ), .D(\mreg/_06216_ ), .Q(\mreg/rf[8][27] ), .QN(\mreg/_05680_ ) );
DFF_X1 \mreg/_11078_ ( .CK(clk ), .D(\mreg/_06217_ ), .Q(\mreg/rf[8][28] ), .QN(\mreg/_05679_ ) );
DFF_X1 \mreg/_11079_ ( .CK(clk ), .D(\mreg/_06218_ ), .Q(\mreg/rf[8][29] ), .QN(\mreg/_05678_ ) );
DFF_X1 \mreg/_11080_ ( .CK(clk ), .D(\mreg/_06219_ ), .Q(\mreg/rf[8][30] ), .QN(\mreg/_05677_ ) );
DFF_X1 \mreg/_11081_ ( .CK(clk ), .D(\mreg/_06220_ ), .Q(\mreg/rf[8][31] ), .QN(\mreg/_05676_ ) );
DFF_X1 \mreg/_11082_ ( .CK(clk ), .D(\mreg/_06221_ ), .Q(\mreg/rf[9][0] ), .QN(\mreg/_05675_ ) );
DFF_X1 \mreg/_11083_ ( .CK(clk ), .D(\mreg/_06222_ ), .Q(\mreg/rf[9][1] ), .QN(\mreg/_05674_ ) );
DFF_X1 \mreg/_11084_ ( .CK(clk ), .D(\mreg/_06223_ ), .Q(\mreg/rf[9][2] ), .QN(\mreg/_05673_ ) );
DFF_X1 \mreg/_11085_ ( .CK(clk ), .D(\mreg/_06224_ ), .Q(\mreg/rf[9][3] ), .QN(\mreg/_05672_ ) );
DFF_X1 \mreg/_11086_ ( .CK(clk ), .D(\mreg/_06225_ ), .Q(\mreg/rf[9][4] ), .QN(\mreg/_05671_ ) );
DFF_X1 \mreg/_11087_ ( .CK(clk ), .D(\mreg/_06226_ ), .Q(\mreg/rf[9][5] ), .QN(\mreg/_05670_ ) );
DFF_X1 \mreg/_11088_ ( .CK(clk ), .D(\mreg/_06227_ ), .Q(\mreg/rf[9][6] ), .QN(\mreg/_05669_ ) );
DFF_X1 \mreg/_11089_ ( .CK(clk ), .D(\mreg/_06228_ ), .Q(\mreg/rf[9][7] ), .QN(\mreg/_05668_ ) );
DFF_X1 \mreg/_11090_ ( .CK(clk ), .D(\mreg/_06229_ ), .Q(\mreg/rf[9][8] ), .QN(\mreg/_05667_ ) );
DFF_X1 \mreg/_11091_ ( .CK(clk ), .D(\mreg/_06230_ ), .Q(\mreg/rf[9][9] ), .QN(\mreg/_05666_ ) );
DFF_X1 \mreg/_11092_ ( .CK(clk ), .D(\mreg/_06231_ ), .Q(\mreg/rf[9][10] ), .QN(\mreg/_05665_ ) );
DFF_X1 \mreg/_11093_ ( .CK(clk ), .D(\mreg/_06232_ ), .Q(\mreg/rf[9][11] ), .QN(\mreg/_05664_ ) );
DFF_X1 \mreg/_11094_ ( .CK(clk ), .D(\mreg/_06233_ ), .Q(\mreg/rf[9][12] ), .QN(\mreg/_05663_ ) );
DFF_X1 \mreg/_11095_ ( .CK(clk ), .D(\mreg/_06234_ ), .Q(\mreg/rf[9][13] ), .QN(\mreg/_05662_ ) );
DFF_X1 \mreg/_11096_ ( .CK(clk ), .D(\mreg/_06235_ ), .Q(\mreg/rf[9][14] ), .QN(\mreg/_05661_ ) );
DFF_X1 \mreg/_11097_ ( .CK(clk ), .D(\mreg/_06236_ ), .Q(\mreg/rf[9][15] ), .QN(\mreg/_05660_ ) );
DFF_X1 \mreg/_11098_ ( .CK(clk ), .D(\mreg/_06237_ ), .Q(\mreg/rf[9][16] ), .QN(\mreg/_05659_ ) );
DFF_X1 \mreg/_11099_ ( .CK(clk ), .D(\mreg/_06238_ ), .Q(\mreg/rf[9][17] ), .QN(\mreg/_05658_ ) );
DFF_X1 \mreg/_11100_ ( .CK(clk ), .D(\mreg/_06239_ ), .Q(\mreg/rf[9][18] ), .QN(\mreg/_05657_ ) );
DFF_X1 \mreg/_11101_ ( .CK(clk ), .D(\mreg/_06240_ ), .Q(\mreg/rf[9][19] ), .QN(\mreg/_05656_ ) );
DFF_X1 \mreg/_11102_ ( .CK(clk ), .D(\mreg/_06241_ ), .Q(\mreg/rf[9][20] ), .QN(\mreg/_05655_ ) );
DFF_X1 \mreg/_11103_ ( .CK(clk ), .D(\mreg/_06242_ ), .Q(\mreg/rf[9][21] ), .QN(\mreg/_05654_ ) );
DFF_X1 \mreg/_11104_ ( .CK(clk ), .D(\mreg/_06243_ ), .Q(\mreg/rf[9][22] ), .QN(\mreg/_05653_ ) );
DFF_X1 \mreg/_11105_ ( .CK(clk ), .D(\mreg/_06244_ ), .Q(\mreg/rf[9][23] ), .QN(\mreg/_05652_ ) );
DFF_X1 \mreg/_11106_ ( .CK(clk ), .D(\mreg/_06245_ ), .Q(\mreg/rf[9][24] ), .QN(\mreg/_05651_ ) );
DFF_X1 \mreg/_11107_ ( .CK(clk ), .D(\mreg/_06246_ ), .Q(\mreg/rf[9][25] ), .QN(\mreg/_05650_ ) );
DFF_X1 \mreg/_11108_ ( .CK(clk ), .D(\mreg/_06247_ ), .Q(\mreg/rf[9][26] ), .QN(\mreg/_05649_ ) );
DFF_X1 \mreg/_11109_ ( .CK(clk ), .D(\mreg/_06248_ ), .Q(\mreg/rf[9][27] ), .QN(\mreg/_05648_ ) );
DFF_X1 \mreg/_11110_ ( .CK(clk ), .D(\mreg/_06249_ ), .Q(\mreg/rf[9][28] ), .QN(\mreg/_05647_ ) );
DFF_X1 \mreg/_11111_ ( .CK(clk ), .D(\mreg/_06250_ ), .Q(\mreg/rf[9][29] ), .QN(\mreg/_05646_ ) );
DFF_X1 \mreg/_11112_ ( .CK(clk ), .D(\mreg/_06251_ ), .Q(\mreg/rf[9][30] ), .QN(\mreg/_05645_ ) );
DFF_X1 \mreg/_11113_ ( .CK(clk ), .D(\mreg/_06252_ ), .Q(\mreg/rf[9][31] ), .QN(\mreg/_05644_ ) );
DFF_X1 \mreg/_11114_ ( .CK(clk ), .D(\mreg/_06253_ ), .Q(\mreg/rf[10][0] ), .QN(\mreg/_05643_ ) );
DFF_X1 \mreg/_11115_ ( .CK(clk ), .D(\mreg/_06254_ ), .Q(\mreg/rf[10][1] ), .QN(\mreg/_05642_ ) );
DFF_X1 \mreg/_11116_ ( .CK(clk ), .D(\mreg/_06255_ ), .Q(\mreg/rf[10][2] ), .QN(\mreg/_05641_ ) );
DFF_X1 \mreg/_11117_ ( .CK(clk ), .D(\mreg/_06256_ ), .Q(\mreg/rf[10][3] ), .QN(\mreg/_05640_ ) );
DFF_X1 \mreg/_11118_ ( .CK(clk ), .D(\mreg/_06257_ ), .Q(\mreg/rf[10][4] ), .QN(\mreg/_05639_ ) );
DFF_X1 \mreg/_11119_ ( .CK(clk ), .D(\mreg/_06258_ ), .Q(\mreg/rf[10][5] ), .QN(\mreg/_05638_ ) );
DFF_X1 \mreg/_11120_ ( .CK(clk ), .D(\mreg/_06259_ ), .Q(\mreg/rf[10][6] ), .QN(\mreg/_05637_ ) );
DFF_X1 \mreg/_11121_ ( .CK(clk ), .D(\mreg/_06260_ ), .Q(\mreg/rf[10][7] ), .QN(\mreg/_05636_ ) );
DFF_X1 \mreg/_11122_ ( .CK(clk ), .D(\mreg/_06261_ ), .Q(\mreg/rf[10][8] ), .QN(\mreg/_05635_ ) );
DFF_X1 \mreg/_11123_ ( .CK(clk ), .D(\mreg/_06262_ ), .Q(\mreg/rf[10][9] ), .QN(\mreg/_05634_ ) );
DFF_X1 \mreg/_11124_ ( .CK(clk ), .D(\mreg/_06263_ ), .Q(\mreg/rf[10][10] ), .QN(\mreg/_05633_ ) );
DFF_X1 \mreg/_11125_ ( .CK(clk ), .D(\mreg/_06264_ ), .Q(\mreg/rf[10][11] ), .QN(\mreg/_05632_ ) );
DFF_X1 \mreg/_11126_ ( .CK(clk ), .D(\mreg/_06265_ ), .Q(\mreg/rf[10][12] ), .QN(\mreg/_05631_ ) );
DFF_X1 \mreg/_11127_ ( .CK(clk ), .D(\mreg/_06266_ ), .Q(\mreg/rf[10][13] ), .QN(\mreg/_05630_ ) );
DFF_X1 \mreg/_11128_ ( .CK(clk ), .D(\mreg/_06267_ ), .Q(\mreg/rf[10][14] ), .QN(\mreg/_05629_ ) );
DFF_X1 \mreg/_11129_ ( .CK(clk ), .D(\mreg/_06268_ ), .Q(\mreg/rf[10][15] ), .QN(\mreg/_05628_ ) );
DFF_X1 \mreg/_11130_ ( .CK(clk ), .D(\mreg/_06269_ ), .Q(\mreg/rf[10][16] ), .QN(\mreg/_05627_ ) );
DFF_X1 \mreg/_11131_ ( .CK(clk ), .D(\mreg/_06270_ ), .Q(\mreg/rf[10][17] ), .QN(\mreg/_05626_ ) );
DFF_X1 \mreg/_11132_ ( .CK(clk ), .D(\mreg/_06271_ ), .Q(\mreg/rf[10][18] ), .QN(\mreg/_05625_ ) );
DFF_X1 \mreg/_11133_ ( .CK(clk ), .D(\mreg/_06272_ ), .Q(\mreg/rf[10][19] ), .QN(\mreg/_05624_ ) );
DFF_X1 \mreg/_11134_ ( .CK(clk ), .D(\mreg/_06273_ ), .Q(\mreg/rf[10][20] ), .QN(\mreg/_05623_ ) );
DFF_X1 \mreg/_11135_ ( .CK(clk ), .D(\mreg/_06274_ ), .Q(\mreg/rf[10][21] ), .QN(\mreg/_05622_ ) );
DFF_X1 \mreg/_11136_ ( .CK(clk ), .D(\mreg/_06275_ ), .Q(\mreg/rf[10][22] ), .QN(\mreg/_05621_ ) );
DFF_X1 \mreg/_11137_ ( .CK(clk ), .D(\mreg/_06276_ ), .Q(\mreg/rf[10][23] ), .QN(\mreg/_05620_ ) );
DFF_X1 \mreg/_11138_ ( .CK(clk ), .D(\mreg/_06277_ ), .Q(\mreg/rf[10][24] ), .QN(\mreg/_05619_ ) );
DFF_X1 \mreg/_11139_ ( .CK(clk ), .D(\mreg/_06278_ ), .Q(\mreg/rf[10][25] ), .QN(\mreg/_05618_ ) );
DFF_X1 \mreg/_11140_ ( .CK(clk ), .D(\mreg/_06279_ ), .Q(\mreg/rf[10][26] ), .QN(\mreg/_05617_ ) );
DFF_X1 \mreg/_11141_ ( .CK(clk ), .D(\mreg/_06280_ ), .Q(\mreg/rf[10][27] ), .QN(\mreg/_05616_ ) );
DFF_X1 \mreg/_11142_ ( .CK(clk ), .D(\mreg/_06281_ ), .Q(\mreg/rf[10][28] ), .QN(\mreg/_05615_ ) );
DFF_X1 \mreg/_11143_ ( .CK(clk ), .D(\mreg/_06282_ ), .Q(\mreg/rf[10][29] ), .QN(\mreg/_05614_ ) );
DFF_X1 \mreg/_11144_ ( .CK(clk ), .D(\mreg/_06283_ ), .Q(\mreg/rf[10][30] ), .QN(\mreg/_05613_ ) );
DFF_X1 \mreg/_11145_ ( .CK(clk ), .D(\mreg/_06284_ ), .Q(\mreg/rf[10][31] ), .QN(\mreg/_05612_ ) );
DFF_X1 \mreg/_11146_ ( .CK(clk ), .D(\mreg/_06285_ ), .Q(\mreg/rf[11][0] ), .QN(\mreg/_05611_ ) );
DFF_X1 \mreg/_11147_ ( .CK(clk ), .D(\mreg/_06286_ ), .Q(\mreg/rf[11][1] ), .QN(\mreg/_05610_ ) );
DFF_X1 \mreg/_11148_ ( .CK(clk ), .D(\mreg/_06287_ ), .Q(\mreg/rf[11][2] ), .QN(\mreg/_05609_ ) );
DFF_X1 \mreg/_11149_ ( .CK(clk ), .D(\mreg/_06288_ ), .Q(\mreg/rf[11][3] ), .QN(\mreg/_05608_ ) );
DFF_X1 \mreg/_11150_ ( .CK(clk ), .D(\mreg/_06289_ ), .Q(\mreg/rf[11][4] ), .QN(\mreg/_05607_ ) );
DFF_X1 \mreg/_11151_ ( .CK(clk ), .D(\mreg/_06290_ ), .Q(\mreg/rf[11][5] ), .QN(\mreg/_05606_ ) );
DFF_X1 \mreg/_11152_ ( .CK(clk ), .D(\mreg/_06291_ ), .Q(\mreg/rf[11][6] ), .QN(\mreg/_05605_ ) );
DFF_X1 \mreg/_11153_ ( .CK(clk ), .D(\mreg/_06292_ ), .Q(\mreg/rf[11][7] ), .QN(\mreg/_05604_ ) );
DFF_X1 \mreg/_11154_ ( .CK(clk ), .D(\mreg/_06293_ ), .Q(\mreg/rf[11][8] ), .QN(\mreg/_05603_ ) );
DFF_X1 \mreg/_11155_ ( .CK(clk ), .D(\mreg/_06294_ ), .Q(\mreg/rf[11][9] ), .QN(\mreg/_05602_ ) );
DFF_X1 \mreg/_11156_ ( .CK(clk ), .D(\mreg/_06295_ ), .Q(\mreg/rf[11][10] ), .QN(\mreg/_05601_ ) );
DFF_X1 \mreg/_11157_ ( .CK(clk ), .D(\mreg/_06296_ ), .Q(\mreg/rf[11][11] ), .QN(\mreg/_05600_ ) );
DFF_X1 \mreg/_11158_ ( .CK(clk ), .D(\mreg/_06297_ ), .Q(\mreg/rf[11][12] ), .QN(\mreg/_05599_ ) );
DFF_X1 \mreg/_11159_ ( .CK(clk ), .D(\mreg/_06298_ ), .Q(\mreg/rf[11][13] ), .QN(\mreg/_05598_ ) );
DFF_X1 \mreg/_11160_ ( .CK(clk ), .D(\mreg/_06299_ ), .Q(\mreg/rf[11][14] ), .QN(\mreg/_05597_ ) );
DFF_X1 \mreg/_11161_ ( .CK(clk ), .D(\mreg/_06300_ ), .Q(\mreg/rf[11][15] ), .QN(\mreg/_05596_ ) );
DFF_X1 \mreg/_11162_ ( .CK(clk ), .D(\mreg/_06301_ ), .Q(\mreg/rf[11][16] ), .QN(\mreg/_05595_ ) );
DFF_X1 \mreg/_11163_ ( .CK(clk ), .D(\mreg/_06302_ ), .Q(\mreg/rf[11][17] ), .QN(\mreg/_05594_ ) );
DFF_X1 \mreg/_11164_ ( .CK(clk ), .D(\mreg/_06303_ ), .Q(\mreg/rf[11][18] ), .QN(\mreg/_05593_ ) );
DFF_X1 \mreg/_11165_ ( .CK(clk ), .D(\mreg/_06304_ ), .Q(\mreg/rf[11][19] ), .QN(\mreg/_05592_ ) );
DFF_X1 \mreg/_11166_ ( .CK(clk ), .D(\mreg/_06305_ ), .Q(\mreg/rf[11][20] ), .QN(\mreg/_05591_ ) );
DFF_X1 \mreg/_11167_ ( .CK(clk ), .D(\mreg/_06306_ ), .Q(\mreg/rf[11][21] ), .QN(\mreg/_05590_ ) );
DFF_X1 \mreg/_11168_ ( .CK(clk ), .D(\mreg/_06307_ ), .Q(\mreg/rf[11][22] ), .QN(\mreg/_05589_ ) );
DFF_X1 \mreg/_11169_ ( .CK(clk ), .D(\mreg/_06308_ ), .Q(\mreg/rf[11][23] ), .QN(\mreg/_05588_ ) );
DFF_X1 \mreg/_11170_ ( .CK(clk ), .D(\mreg/_06309_ ), .Q(\mreg/rf[11][24] ), .QN(\mreg/_05587_ ) );
DFF_X1 \mreg/_11171_ ( .CK(clk ), .D(\mreg/_06310_ ), .Q(\mreg/rf[11][25] ), .QN(\mreg/_05586_ ) );
DFF_X1 \mreg/_11172_ ( .CK(clk ), .D(\mreg/_06311_ ), .Q(\mreg/rf[11][26] ), .QN(\mreg/_05585_ ) );
DFF_X1 \mreg/_11173_ ( .CK(clk ), .D(\mreg/_06312_ ), .Q(\mreg/rf[11][27] ), .QN(\mreg/_05584_ ) );
DFF_X1 \mreg/_11174_ ( .CK(clk ), .D(\mreg/_06313_ ), .Q(\mreg/rf[11][28] ), .QN(\mreg/_05583_ ) );
DFF_X1 \mreg/_11175_ ( .CK(clk ), .D(\mreg/_06314_ ), .Q(\mreg/rf[11][29] ), .QN(\mreg/_05582_ ) );
DFF_X1 \mreg/_11176_ ( .CK(clk ), .D(\mreg/_06315_ ), .Q(\mreg/rf[11][30] ), .QN(\mreg/_05581_ ) );
DFF_X1 \mreg/_11177_ ( .CK(clk ), .D(\mreg/_06316_ ), .Q(\mreg/rf[11][31] ), .QN(\mreg/_05580_ ) );
DFF_X1 \mreg/_11178_ ( .CK(clk ), .D(\mreg/_06317_ ), .Q(\mreg/rf[12][0] ), .QN(\mreg/_05579_ ) );
DFF_X1 \mreg/_11179_ ( .CK(clk ), .D(\mreg/_06318_ ), .Q(\mreg/rf[12][1] ), .QN(\mreg/_05578_ ) );
DFF_X1 \mreg/_11180_ ( .CK(clk ), .D(\mreg/_06319_ ), .Q(\mreg/rf[12][2] ), .QN(\mreg/_05577_ ) );
DFF_X1 \mreg/_11181_ ( .CK(clk ), .D(\mreg/_06320_ ), .Q(\mreg/rf[12][3] ), .QN(\mreg/_05576_ ) );
DFF_X1 \mreg/_11182_ ( .CK(clk ), .D(\mreg/_06321_ ), .Q(\mreg/rf[12][4] ), .QN(\mreg/_05575_ ) );
DFF_X1 \mreg/_11183_ ( .CK(clk ), .D(\mreg/_06322_ ), .Q(\mreg/rf[12][5] ), .QN(\mreg/_05574_ ) );
DFF_X1 \mreg/_11184_ ( .CK(clk ), .D(\mreg/_06323_ ), .Q(\mreg/rf[12][6] ), .QN(\mreg/_05573_ ) );
DFF_X1 \mreg/_11185_ ( .CK(clk ), .D(\mreg/_06324_ ), .Q(\mreg/rf[12][7] ), .QN(\mreg/_05572_ ) );
DFF_X1 \mreg/_11186_ ( .CK(clk ), .D(\mreg/_06325_ ), .Q(\mreg/rf[12][8] ), .QN(\mreg/_05571_ ) );
DFF_X1 \mreg/_11187_ ( .CK(clk ), .D(\mreg/_06326_ ), .Q(\mreg/rf[12][9] ), .QN(\mreg/_05570_ ) );
DFF_X1 \mreg/_11188_ ( .CK(clk ), .D(\mreg/_06327_ ), .Q(\mreg/rf[12][10] ), .QN(\mreg/_05569_ ) );
DFF_X1 \mreg/_11189_ ( .CK(clk ), .D(\mreg/_06328_ ), .Q(\mreg/rf[12][11] ), .QN(\mreg/_05568_ ) );
DFF_X1 \mreg/_11190_ ( .CK(clk ), .D(\mreg/_06329_ ), .Q(\mreg/rf[12][12] ), .QN(\mreg/_05567_ ) );
DFF_X1 \mreg/_11191_ ( .CK(clk ), .D(\mreg/_06330_ ), .Q(\mreg/rf[12][13] ), .QN(\mreg/_05566_ ) );
DFF_X1 \mreg/_11192_ ( .CK(clk ), .D(\mreg/_06331_ ), .Q(\mreg/rf[12][14] ), .QN(\mreg/_05565_ ) );
DFF_X1 \mreg/_11193_ ( .CK(clk ), .D(\mreg/_06332_ ), .Q(\mreg/rf[12][15] ), .QN(\mreg/_05564_ ) );
DFF_X1 \mreg/_11194_ ( .CK(clk ), .D(\mreg/_06333_ ), .Q(\mreg/rf[12][16] ), .QN(\mreg/_05563_ ) );
DFF_X1 \mreg/_11195_ ( .CK(clk ), .D(\mreg/_06334_ ), .Q(\mreg/rf[12][17] ), .QN(\mreg/_05562_ ) );
DFF_X1 \mreg/_11196_ ( .CK(clk ), .D(\mreg/_06335_ ), .Q(\mreg/rf[12][18] ), .QN(\mreg/_05561_ ) );
DFF_X1 \mreg/_11197_ ( .CK(clk ), .D(\mreg/_06336_ ), .Q(\mreg/rf[12][19] ), .QN(\mreg/_05560_ ) );
DFF_X1 \mreg/_11198_ ( .CK(clk ), .D(\mreg/_06337_ ), .Q(\mreg/rf[12][20] ), .QN(\mreg/_05559_ ) );
DFF_X1 \mreg/_11199_ ( .CK(clk ), .D(\mreg/_06338_ ), .Q(\mreg/rf[12][21] ), .QN(\mreg/_05558_ ) );
DFF_X1 \mreg/_11200_ ( .CK(clk ), .D(\mreg/_06339_ ), .Q(\mreg/rf[12][22] ), .QN(\mreg/_05557_ ) );
DFF_X1 \mreg/_11201_ ( .CK(clk ), .D(\mreg/_06340_ ), .Q(\mreg/rf[12][23] ), .QN(\mreg/_05556_ ) );
DFF_X1 \mreg/_11202_ ( .CK(clk ), .D(\mreg/_06341_ ), .Q(\mreg/rf[12][24] ), .QN(\mreg/_05555_ ) );
DFF_X1 \mreg/_11203_ ( .CK(clk ), .D(\mreg/_06342_ ), .Q(\mreg/rf[12][25] ), .QN(\mreg/_05554_ ) );
DFF_X1 \mreg/_11204_ ( .CK(clk ), .D(\mreg/_06343_ ), .Q(\mreg/rf[12][26] ), .QN(\mreg/_05553_ ) );
DFF_X1 \mreg/_11205_ ( .CK(clk ), .D(\mreg/_06344_ ), .Q(\mreg/rf[12][27] ), .QN(\mreg/_05552_ ) );
DFF_X1 \mreg/_11206_ ( .CK(clk ), .D(\mreg/_06345_ ), .Q(\mreg/rf[12][28] ), .QN(\mreg/_05551_ ) );
DFF_X1 \mreg/_11207_ ( .CK(clk ), .D(\mreg/_06346_ ), .Q(\mreg/rf[12][29] ), .QN(\mreg/_05550_ ) );
DFF_X1 \mreg/_11208_ ( .CK(clk ), .D(\mreg/_06347_ ), .Q(\mreg/rf[12][30] ), .QN(\mreg/_05549_ ) );
DFF_X1 \mreg/_11209_ ( .CK(clk ), .D(\mreg/_06348_ ), .Q(\mreg/rf[12][31] ), .QN(\mreg/_05548_ ) );
DFF_X1 \mreg/_11210_ ( .CK(clk ), .D(\mreg/_06349_ ), .Q(\mreg/rf[13][0] ), .QN(\mreg/_05547_ ) );
DFF_X1 \mreg/_11211_ ( .CK(clk ), .D(\mreg/_06350_ ), .Q(\mreg/rf[13][1] ), .QN(\mreg/_05546_ ) );
DFF_X1 \mreg/_11212_ ( .CK(clk ), .D(\mreg/_06351_ ), .Q(\mreg/rf[13][2] ), .QN(\mreg/_05545_ ) );
DFF_X1 \mreg/_11213_ ( .CK(clk ), .D(\mreg/_06352_ ), .Q(\mreg/rf[13][3] ), .QN(\mreg/_05544_ ) );
DFF_X1 \mreg/_11214_ ( .CK(clk ), .D(\mreg/_06353_ ), .Q(\mreg/rf[13][4] ), .QN(\mreg/_05543_ ) );
DFF_X1 \mreg/_11215_ ( .CK(clk ), .D(\mreg/_06354_ ), .Q(\mreg/rf[13][5] ), .QN(\mreg/_05542_ ) );
DFF_X1 \mreg/_11216_ ( .CK(clk ), .D(\mreg/_06355_ ), .Q(\mreg/rf[13][6] ), .QN(\mreg/_05541_ ) );
DFF_X1 \mreg/_11217_ ( .CK(clk ), .D(\mreg/_06356_ ), .Q(\mreg/rf[13][7] ), .QN(\mreg/_05540_ ) );
DFF_X1 \mreg/_11218_ ( .CK(clk ), .D(\mreg/_06357_ ), .Q(\mreg/rf[13][8] ), .QN(\mreg/_05539_ ) );
DFF_X1 \mreg/_11219_ ( .CK(clk ), .D(\mreg/_06358_ ), .Q(\mreg/rf[13][9] ), .QN(\mreg/_05538_ ) );
DFF_X1 \mreg/_11220_ ( .CK(clk ), .D(\mreg/_06359_ ), .Q(\mreg/rf[13][10] ), .QN(\mreg/_05537_ ) );
DFF_X1 \mreg/_11221_ ( .CK(clk ), .D(\mreg/_06360_ ), .Q(\mreg/rf[13][11] ), .QN(\mreg/_05536_ ) );
DFF_X1 \mreg/_11222_ ( .CK(clk ), .D(\mreg/_06361_ ), .Q(\mreg/rf[13][12] ), .QN(\mreg/_05535_ ) );
DFF_X1 \mreg/_11223_ ( .CK(clk ), .D(\mreg/_06362_ ), .Q(\mreg/rf[13][13] ), .QN(\mreg/_05534_ ) );
DFF_X1 \mreg/_11224_ ( .CK(clk ), .D(\mreg/_06363_ ), .Q(\mreg/rf[13][14] ), .QN(\mreg/_05533_ ) );
DFF_X1 \mreg/_11225_ ( .CK(clk ), .D(\mreg/_06364_ ), .Q(\mreg/rf[13][15] ), .QN(\mreg/_05532_ ) );
DFF_X1 \mreg/_11226_ ( .CK(clk ), .D(\mreg/_06365_ ), .Q(\mreg/rf[13][16] ), .QN(\mreg/_05531_ ) );
DFF_X1 \mreg/_11227_ ( .CK(clk ), .D(\mreg/_06366_ ), .Q(\mreg/rf[13][17] ), .QN(\mreg/_05530_ ) );
DFF_X1 \mreg/_11228_ ( .CK(clk ), .D(\mreg/_06367_ ), .Q(\mreg/rf[13][18] ), .QN(\mreg/_05529_ ) );
DFF_X1 \mreg/_11229_ ( .CK(clk ), .D(\mreg/_06368_ ), .Q(\mreg/rf[13][19] ), .QN(\mreg/_05528_ ) );
DFF_X1 \mreg/_11230_ ( .CK(clk ), .D(\mreg/_06369_ ), .Q(\mreg/rf[13][20] ), .QN(\mreg/_05527_ ) );
DFF_X1 \mreg/_11231_ ( .CK(clk ), .D(\mreg/_06370_ ), .Q(\mreg/rf[13][21] ), .QN(\mreg/_05526_ ) );
DFF_X1 \mreg/_11232_ ( .CK(clk ), .D(\mreg/_06371_ ), .Q(\mreg/rf[13][22] ), .QN(\mreg/_05525_ ) );
DFF_X1 \mreg/_11233_ ( .CK(clk ), .D(\mreg/_06372_ ), .Q(\mreg/rf[13][23] ), .QN(\mreg/_05524_ ) );
DFF_X1 \mreg/_11234_ ( .CK(clk ), .D(\mreg/_06373_ ), .Q(\mreg/rf[13][24] ), .QN(\mreg/_05523_ ) );
DFF_X1 \mreg/_11235_ ( .CK(clk ), .D(\mreg/_06374_ ), .Q(\mreg/rf[13][25] ), .QN(\mreg/_05522_ ) );
DFF_X1 \mreg/_11236_ ( .CK(clk ), .D(\mreg/_06375_ ), .Q(\mreg/rf[13][26] ), .QN(\mreg/_05521_ ) );
DFF_X1 \mreg/_11237_ ( .CK(clk ), .D(\mreg/_06376_ ), .Q(\mreg/rf[13][27] ), .QN(\mreg/_05520_ ) );
DFF_X1 \mreg/_11238_ ( .CK(clk ), .D(\mreg/_06377_ ), .Q(\mreg/rf[13][28] ), .QN(\mreg/_05519_ ) );
DFF_X1 \mreg/_11239_ ( .CK(clk ), .D(\mreg/_06378_ ), .Q(\mreg/rf[13][29] ), .QN(\mreg/_05518_ ) );
DFF_X1 \mreg/_11240_ ( .CK(clk ), .D(\mreg/_06379_ ), .Q(\mreg/rf[13][30] ), .QN(\mreg/_05517_ ) );
DFF_X1 \mreg/_11241_ ( .CK(clk ), .D(\mreg/_06380_ ), .Q(\mreg/rf[13][31] ), .QN(\mreg/_05516_ ) );
DFF_X1 \mreg/_11242_ ( .CK(clk ), .D(\mreg/_06381_ ), .Q(\mreg/rf[14][0] ), .QN(\mreg/_05515_ ) );
DFF_X1 \mreg/_11243_ ( .CK(clk ), .D(\mreg/_06382_ ), .Q(\mreg/rf[14][1] ), .QN(\mreg/_05514_ ) );
DFF_X1 \mreg/_11244_ ( .CK(clk ), .D(\mreg/_06383_ ), .Q(\mreg/rf[14][2] ), .QN(\mreg/_05513_ ) );
DFF_X1 \mreg/_11245_ ( .CK(clk ), .D(\mreg/_06384_ ), .Q(\mreg/rf[14][3] ), .QN(\mreg/_05512_ ) );
DFF_X1 \mreg/_11246_ ( .CK(clk ), .D(\mreg/_06385_ ), .Q(\mreg/rf[14][4] ), .QN(\mreg/_05511_ ) );
DFF_X1 \mreg/_11247_ ( .CK(clk ), .D(\mreg/_06386_ ), .Q(\mreg/rf[14][5] ), .QN(\mreg/_05510_ ) );
DFF_X1 \mreg/_11248_ ( .CK(clk ), .D(\mreg/_06387_ ), .Q(\mreg/rf[14][6] ), .QN(\mreg/_05509_ ) );
DFF_X1 \mreg/_11249_ ( .CK(clk ), .D(\mreg/_06388_ ), .Q(\mreg/rf[14][7] ), .QN(\mreg/_05508_ ) );
DFF_X1 \mreg/_11250_ ( .CK(clk ), .D(\mreg/_06389_ ), .Q(\mreg/rf[14][8] ), .QN(\mreg/_05507_ ) );
DFF_X1 \mreg/_11251_ ( .CK(clk ), .D(\mreg/_06390_ ), .Q(\mreg/rf[14][9] ), .QN(\mreg/_05506_ ) );
DFF_X1 \mreg/_11252_ ( .CK(clk ), .D(\mreg/_06391_ ), .Q(\mreg/rf[14][10] ), .QN(\mreg/_05505_ ) );
DFF_X1 \mreg/_11253_ ( .CK(clk ), .D(\mreg/_06392_ ), .Q(\mreg/rf[14][11] ), .QN(\mreg/_05504_ ) );
DFF_X1 \mreg/_11254_ ( .CK(clk ), .D(\mreg/_06393_ ), .Q(\mreg/rf[14][12] ), .QN(\mreg/_05503_ ) );
DFF_X1 \mreg/_11255_ ( .CK(clk ), .D(\mreg/_06394_ ), .Q(\mreg/rf[14][13] ), .QN(\mreg/_05502_ ) );
DFF_X1 \mreg/_11256_ ( .CK(clk ), .D(\mreg/_06395_ ), .Q(\mreg/rf[14][14] ), .QN(\mreg/_05501_ ) );
DFF_X1 \mreg/_11257_ ( .CK(clk ), .D(\mreg/_06396_ ), .Q(\mreg/rf[14][15] ), .QN(\mreg/_05500_ ) );
DFF_X1 \mreg/_11258_ ( .CK(clk ), .D(\mreg/_06397_ ), .Q(\mreg/rf[14][16] ), .QN(\mreg/_05499_ ) );
DFF_X1 \mreg/_11259_ ( .CK(clk ), .D(\mreg/_06398_ ), .Q(\mreg/rf[14][17] ), .QN(\mreg/_05498_ ) );
DFF_X1 \mreg/_11260_ ( .CK(clk ), .D(\mreg/_06399_ ), .Q(\mreg/rf[14][18] ), .QN(\mreg/_05497_ ) );
DFF_X1 \mreg/_11261_ ( .CK(clk ), .D(\mreg/_06400_ ), .Q(\mreg/rf[14][19] ), .QN(\mreg/_05496_ ) );
DFF_X1 \mreg/_11262_ ( .CK(clk ), .D(\mreg/_06401_ ), .Q(\mreg/rf[14][20] ), .QN(\mreg/_05495_ ) );
DFF_X1 \mreg/_11263_ ( .CK(clk ), .D(\mreg/_06402_ ), .Q(\mreg/rf[14][21] ), .QN(\mreg/_05494_ ) );
DFF_X1 \mreg/_11264_ ( .CK(clk ), .D(\mreg/_06403_ ), .Q(\mreg/rf[14][22] ), .QN(\mreg/_05493_ ) );
DFF_X1 \mreg/_11265_ ( .CK(clk ), .D(\mreg/_06404_ ), .Q(\mreg/rf[14][23] ), .QN(\mreg/_05492_ ) );
DFF_X1 \mreg/_11266_ ( .CK(clk ), .D(\mreg/_06405_ ), .Q(\mreg/rf[14][24] ), .QN(\mreg/_05491_ ) );
DFF_X1 \mreg/_11267_ ( .CK(clk ), .D(\mreg/_06406_ ), .Q(\mreg/rf[14][25] ), .QN(\mreg/_05490_ ) );
DFF_X1 \mreg/_11268_ ( .CK(clk ), .D(\mreg/_06407_ ), .Q(\mreg/rf[14][26] ), .QN(\mreg/_05489_ ) );
DFF_X1 \mreg/_11269_ ( .CK(clk ), .D(\mreg/_06408_ ), .Q(\mreg/rf[14][27] ), .QN(\mreg/_05488_ ) );
DFF_X1 \mreg/_11270_ ( .CK(clk ), .D(\mreg/_06409_ ), .Q(\mreg/rf[14][28] ), .QN(\mreg/_05487_ ) );
DFF_X1 \mreg/_11271_ ( .CK(clk ), .D(\mreg/_06410_ ), .Q(\mreg/rf[14][29] ), .QN(\mreg/_05486_ ) );
DFF_X1 \mreg/_11272_ ( .CK(clk ), .D(\mreg/_06411_ ), .Q(\mreg/rf[14][30] ), .QN(\mreg/_05485_ ) );
DFF_X1 \mreg/_11273_ ( .CK(clk ), .D(\mreg/_06412_ ), .Q(\mreg/rf[14][31] ), .QN(\mreg/_05484_ ) );
DFF_X1 \mreg/_11274_ ( .CK(clk ), .D(\mreg/_06413_ ), .Q(\mreg/rf[15][0] ), .QN(\mreg/_05483_ ) );
DFF_X1 \mreg/_11275_ ( .CK(clk ), .D(\mreg/_06414_ ), .Q(\mreg/rf[15][1] ), .QN(\mreg/_05482_ ) );
DFF_X1 \mreg/_11276_ ( .CK(clk ), .D(\mreg/_06415_ ), .Q(\mreg/rf[15][2] ), .QN(\mreg/_05481_ ) );
DFF_X1 \mreg/_11277_ ( .CK(clk ), .D(\mreg/_06416_ ), .Q(\mreg/rf[15][3] ), .QN(\mreg/_05480_ ) );
DFF_X1 \mreg/_11278_ ( .CK(clk ), .D(\mreg/_06417_ ), .Q(\mreg/rf[15][4] ), .QN(\mreg/_05479_ ) );
DFF_X1 \mreg/_11279_ ( .CK(clk ), .D(\mreg/_06418_ ), .Q(\mreg/rf[15][5] ), .QN(\mreg/_05478_ ) );
DFF_X1 \mreg/_11280_ ( .CK(clk ), .D(\mreg/_06419_ ), .Q(\mreg/rf[15][6] ), .QN(\mreg/_05477_ ) );
DFF_X1 \mreg/_11281_ ( .CK(clk ), .D(\mreg/_06420_ ), .Q(\mreg/rf[15][7] ), .QN(\mreg/_05476_ ) );
DFF_X1 \mreg/_11282_ ( .CK(clk ), .D(\mreg/_06421_ ), .Q(\mreg/rf[15][8] ), .QN(\mreg/_05475_ ) );
DFF_X1 \mreg/_11283_ ( .CK(clk ), .D(\mreg/_06422_ ), .Q(\mreg/rf[15][9] ), .QN(\mreg/_05474_ ) );
DFF_X1 \mreg/_11284_ ( .CK(clk ), .D(\mreg/_06423_ ), .Q(\mreg/rf[15][10] ), .QN(\mreg/_05473_ ) );
DFF_X1 \mreg/_11285_ ( .CK(clk ), .D(\mreg/_06424_ ), .Q(\mreg/rf[15][11] ), .QN(\mreg/_05472_ ) );
DFF_X1 \mreg/_11286_ ( .CK(clk ), .D(\mreg/_06425_ ), .Q(\mreg/rf[15][12] ), .QN(\mreg/_05471_ ) );
DFF_X1 \mreg/_11287_ ( .CK(clk ), .D(\mreg/_06426_ ), .Q(\mreg/rf[15][13] ), .QN(\mreg/_05470_ ) );
DFF_X1 \mreg/_11288_ ( .CK(clk ), .D(\mreg/_06427_ ), .Q(\mreg/rf[15][14] ), .QN(\mreg/_05469_ ) );
DFF_X1 \mreg/_11289_ ( .CK(clk ), .D(\mreg/_06428_ ), .Q(\mreg/rf[15][15] ), .QN(\mreg/_05468_ ) );
DFF_X1 \mreg/_11290_ ( .CK(clk ), .D(\mreg/_06429_ ), .Q(\mreg/rf[15][16] ), .QN(\mreg/_05467_ ) );
DFF_X1 \mreg/_11291_ ( .CK(clk ), .D(\mreg/_06430_ ), .Q(\mreg/rf[15][17] ), .QN(\mreg/_05466_ ) );
DFF_X1 \mreg/_11292_ ( .CK(clk ), .D(\mreg/_06431_ ), .Q(\mreg/rf[15][18] ), .QN(\mreg/_05465_ ) );
DFF_X1 \mreg/_11293_ ( .CK(clk ), .D(\mreg/_06432_ ), .Q(\mreg/rf[15][19] ), .QN(\mreg/_05464_ ) );
DFF_X1 \mreg/_11294_ ( .CK(clk ), .D(\mreg/_06433_ ), .Q(\mreg/rf[15][20] ), .QN(\mreg/_05463_ ) );
DFF_X1 \mreg/_11295_ ( .CK(clk ), .D(\mreg/_06434_ ), .Q(\mreg/rf[15][21] ), .QN(\mreg/_05462_ ) );
DFF_X1 \mreg/_11296_ ( .CK(clk ), .D(\mreg/_06435_ ), .Q(\mreg/rf[15][22] ), .QN(\mreg/_05461_ ) );
DFF_X1 \mreg/_11297_ ( .CK(clk ), .D(\mreg/_06436_ ), .Q(\mreg/rf[15][23] ), .QN(\mreg/_05460_ ) );
DFF_X1 \mreg/_11298_ ( .CK(clk ), .D(\mreg/_06437_ ), .Q(\mreg/rf[15][24] ), .QN(\mreg/_05459_ ) );
DFF_X1 \mreg/_11299_ ( .CK(clk ), .D(\mreg/_06438_ ), .Q(\mreg/rf[15][25] ), .QN(\mreg/_05458_ ) );
DFF_X1 \mreg/_11300_ ( .CK(clk ), .D(\mreg/_06439_ ), .Q(\mreg/rf[15][26] ), .QN(\mreg/_05457_ ) );
DFF_X1 \mreg/_11301_ ( .CK(clk ), .D(\mreg/_06440_ ), .Q(\mreg/rf[15][27] ), .QN(\mreg/_05456_ ) );
DFF_X1 \mreg/_11302_ ( .CK(clk ), .D(\mreg/_06441_ ), .Q(\mreg/rf[15][28] ), .QN(\mreg/_05455_ ) );
DFF_X1 \mreg/_11303_ ( .CK(clk ), .D(\mreg/_06442_ ), .Q(\mreg/rf[15][29] ), .QN(\mreg/_05454_ ) );
DFF_X1 \mreg/_11304_ ( .CK(clk ), .D(\mreg/_06443_ ), .Q(\mreg/rf[15][30] ), .QN(\mreg/_05453_ ) );
DFF_X1 \mreg/_11305_ ( .CK(clk ), .D(\mreg/_06444_ ), .Q(\mreg/rf[15][31] ), .QN(\mreg/_05452_ ) );
DFF_X1 \mreg/_11306_ ( .CK(clk ), .D(\mreg/_06445_ ), .Q(\mreg/rf[16][0] ), .QN(\mreg/_05451_ ) );
DFF_X1 \mreg/_11307_ ( .CK(clk ), .D(\mreg/_06446_ ), .Q(\mreg/rf[16][1] ), .QN(\mreg/_05450_ ) );
DFF_X1 \mreg/_11308_ ( .CK(clk ), .D(\mreg/_06447_ ), .Q(\mreg/rf[16][2] ), .QN(\mreg/_05449_ ) );
DFF_X1 \mreg/_11309_ ( .CK(clk ), .D(\mreg/_06448_ ), .Q(\mreg/rf[16][3] ), .QN(\mreg/_05448_ ) );
DFF_X1 \mreg/_11310_ ( .CK(clk ), .D(\mreg/_06449_ ), .Q(\mreg/rf[16][4] ), .QN(\mreg/_05447_ ) );
DFF_X1 \mreg/_11311_ ( .CK(clk ), .D(\mreg/_06450_ ), .Q(\mreg/rf[16][5] ), .QN(\mreg/_05446_ ) );
DFF_X1 \mreg/_11312_ ( .CK(clk ), .D(\mreg/_06451_ ), .Q(\mreg/rf[16][6] ), .QN(\mreg/_05445_ ) );
DFF_X1 \mreg/_11313_ ( .CK(clk ), .D(\mreg/_06452_ ), .Q(\mreg/rf[16][7] ), .QN(\mreg/_05444_ ) );
DFF_X1 \mreg/_11314_ ( .CK(clk ), .D(\mreg/_06453_ ), .Q(\mreg/rf[16][8] ), .QN(\mreg/_05443_ ) );
DFF_X1 \mreg/_11315_ ( .CK(clk ), .D(\mreg/_06454_ ), .Q(\mreg/rf[16][9] ), .QN(\mreg/_05442_ ) );
DFF_X1 \mreg/_11316_ ( .CK(clk ), .D(\mreg/_06455_ ), .Q(\mreg/rf[16][10] ), .QN(\mreg/_05441_ ) );
DFF_X1 \mreg/_11317_ ( .CK(clk ), .D(\mreg/_06456_ ), .Q(\mreg/rf[16][11] ), .QN(\mreg/_05440_ ) );
DFF_X1 \mreg/_11318_ ( .CK(clk ), .D(\mreg/_06457_ ), .Q(\mreg/rf[16][12] ), .QN(\mreg/_05439_ ) );
DFF_X1 \mreg/_11319_ ( .CK(clk ), .D(\mreg/_06458_ ), .Q(\mreg/rf[16][13] ), .QN(\mreg/_05438_ ) );
DFF_X1 \mreg/_11320_ ( .CK(clk ), .D(\mreg/_06459_ ), .Q(\mreg/rf[16][14] ), .QN(\mreg/_05437_ ) );
DFF_X1 \mreg/_11321_ ( .CK(clk ), .D(\mreg/_06460_ ), .Q(\mreg/rf[16][15] ), .QN(\mreg/_05436_ ) );
DFF_X1 \mreg/_11322_ ( .CK(clk ), .D(\mreg/_06461_ ), .Q(\mreg/rf[16][16] ), .QN(\mreg/_05435_ ) );
DFF_X1 \mreg/_11323_ ( .CK(clk ), .D(\mreg/_06462_ ), .Q(\mreg/rf[16][17] ), .QN(\mreg/_05434_ ) );
DFF_X1 \mreg/_11324_ ( .CK(clk ), .D(\mreg/_06463_ ), .Q(\mreg/rf[16][18] ), .QN(\mreg/_05433_ ) );
DFF_X1 \mreg/_11325_ ( .CK(clk ), .D(\mreg/_06464_ ), .Q(\mreg/rf[16][19] ), .QN(\mreg/_05432_ ) );
DFF_X1 \mreg/_11326_ ( .CK(clk ), .D(\mreg/_06465_ ), .Q(\mreg/rf[16][20] ), .QN(\mreg/_05431_ ) );
DFF_X1 \mreg/_11327_ ( .CK(clk ), .D(\mreg/_06466_ ), .Q(\mreg/rf[16][21] ), .QN(\mreg/_05430_ ) );
DFF_X1 \mreg/_11328_ ( .CK(clk ), .D(\mreg/_06467_ ), .Q(\mreg/rf[16][22] ), .QN(\mreg/_05429_ ) );
DFF_X1 \mreg/_11329_ ( .CK(clk ), .D(\mreg/_06468_ ), .Q(\mreg/rf[16][23] ), .QN(\mreg/_05428_ ) );
DFF_X1 \mreg/_11330_ ( .CK(clk ), .D(\mreg/_06469_ ), .Q(\mreg/rf[16][24] ), .QN(\mreg/_05427_ ) );
DFF_X1 \mreg/_11331_ ( .CK(clk ), .D(\mreg/_06470_ ), .Q(\mreg/rf[16][25] ), .QN(\mreg/_05426_ ) );
DFF_X1 \mreg/_11332_ ( .CK(clk ), .D(\mreg/_06471_ ), .Q(\mreg/rf[16][26] ), .QN(\mreg/_05425_ ) );
DFF_X1 \mreg/_11333_ ( .CK(clk ), .D(\mreg/_06472_ ), .Q(\mreg/rf[16][27] ), .QN(\mreg/_05424_ ) );
DFF_X1 \mreg/_11334_ ( .CK(clk ), .D(\mreg/_06473_ ), .Q(\mreg/rf[16][28] ), .QN(\mreg/_05423_ ) );
DFF_X1 \mreg/_11335_ ( .CK(clk ), .D(\mreg/_06474_ ), .Q(\mreg/rf[16][29] ), .QN(\mreg/_05422_ ) );
DFF_X1 \mreg/_11336_ ( .CK(clk ), .D(\mreg/_06475_ ), .Q(\mreg/rf[16][30] ), .QN(\mreg/_05421_ ) );
DFF_X1 \mreg/_11337_ ( .CK(clk ), .D(\mreg/_06476_ ), .Q(\mreg/rf[16][31] ), .QN(\mreg/_05420_ ) );
DFF_X1 \mreg/_11338_ ( .CK(clk ), .D(\mreg/_06477_ ), .Q(\mreg/rf[17][0] ), .QN(\mreg/_05419_ ) );
DFF_X1 \mreg/_11339_ ( .CK(clk ), .D(\mreg/_06478_ ), .Q(\mreg/rf[17][1] ), .QN(\mreg/_05418_ ) );
DFF_X1 \mreg/_11340_ ( .CK(clk ), .D(\mreg/_06479_ ), .Q(\mreg/rf[17][2] ), .QN(\mreg/_05417_ ) );
DFF_X1 \mreg/_11341_ ( .CK(clk ), .D(\mreg/_06480_ ), .Q(\mreg/rf[17][3] ), .QN(\mreg/_05416_ ) );
DFF_X1 \mreg/_11342_ ( .CK(clk ), .D(\mreg/_06481_ ), .Q(\mreg/rf[17][4] ), .QN(\mreg/_05415_ ) );
DFF_X1 \mreg/_11343_ ( .CK(clk ), .D(\mreg/_06482_ ), .Q(\mreg/rf[17][5] ), .QN(\mreg/_05414_ ) );
DFF_X1 \mreg/_11344_ ( .CK(clk ), .D(\mreg/_06483_ ), .Q(\mreg/rf[17][6] ), .QN(\mreg/_05413_ ) );
DFF_X1 \mreg/_11345_ ( .CK(clk ), .D(\mreg/_06484_ ), .Q(\mreg/rf[17][7] ), .QN(\mreg/_05412_ ) );
DFF_X1 \mreg/_11346_ ( .CK(clk ), .D(\mreg/_06485_ ), .Q(\mreg/rf[17][8] ), .QN(\mreg/_05411_ ) );
DFF_X1 \mreg/_11347_ ( .CK(clk ), .D(\mreg/_06486_ ), .Q(\mreg/rf[17][9] ), .QN(\mreg/_05410_ ) );
DFF_X1 \mreg/_11348_ ( .CK(clk ), .D(\mreg/_06487_ ), .Q(\mreg/rf[17][10] ), .QN(\mreg/_05409_ ) );
DFF_X1 \mreg/_11349_ ( .CK(clk ), .D(\mreg/_06488_ ), .Q(\mreg/rf[17][11] ), .QN(\mreg/_05408_ ) );
DFF_X1 \mreg/_11350_ ( .CK(clk ), .D(\mreg/_06489_ ), .Q(\mreg/rf[17][12] ), .QN(\mreg/_05407_ ) );
DFF_X1 \mreg/_11351_ ( .CK(clk ), .D(\mreg/_06490_ ), .Q(\mreg/rf[17][13] ), .QN(\mreg/_05406_ ) );
DFF_X1 \mreg/_11352_ ( .CK(clk ), .D(\mreg/_06491_ ), .Q(\mreg/rf[17][14] ), .QN(\mreg/_05405_ ) );
DFF_X1 \mreg/_11353_ ( .CK(clk ), .D(\mreg/_06492_ ), .Q(\mreg/rf[17][15] ), .QN(\mreg/_05404_ ) );
DFF_X1 \mreg/_11354_ ( .CK(clk ), .D(\mreg/_06493_ ), .Q(\mreg/rf[17][16] ), .QN(\mreg/_05403_ ) );
DFF_X1 \mreg/_11355_ ( .CK(clk ), .D(\mreg/_06494_ ), .Q(\mreg/rf[17][17] ), .QN(\mreg/_05402_ ) );
DFF_X1 \mreg/_11356_ ( .CK(clk ), .D(\mreg/_06495_ ), .Q(\mreg/rf[17][18] ), .QN(\mreg/_05401_ ) );
DFF_X1 \mreg/_11357_ ( .CK(clk ), .D(\mreg/_06496_ ), .Q(\mreg/rf[17][19] ), .QN(\mreg/_05400_ ) );
DFF_X1 \mreg/_11358_ ( .CK(clk ), .D(\mreg/_06497_ ), .Q(\mreg/rf[17][20] ), .QN(\mreg/_05399_ ) );
DFF_X1 \mreg/_11359_ ( .CK(clk ), .D(\mreg/_06498_ ), .Q(\mreg/rf[17][21] ), .QN(\mreg/_05398_ ) );
DFF_X1 \mreg/_11360_ ( .CK(clk ), .D(\mreg/_06499_ ), .Q(\mreg/rf[17][22] ), .QN(\mreg/_05397_ ) );
DFF_X1 \mreg/_11361_ ( .CK(clk ), .D(\mreg/_06500_ ), .Q(\mreg/rf[17][23] ), .QN(\mreg/_05396_ ) );
DFF_X1 \mreg/_11362_ ( .CK(clk ), .D(\mreg/_06501_ ), .Q(\mreg/rf[17][24] ), .QN(\mreg/_05395_ ) );
DFF_X1 \mreg/_11363_ ( .CK(clk ), .D(\mreg/_06502_ ), .Q(\mreg/rf[17][25] ), .QN(\mreg/_05394_ ) );
DFF_X1 \mreg/_11364_ ( .CK(clk ), .D(\mreg/_06503_ ), .Q(\mreg/rf[17][26] ), .QN(\mreg/_05393_ ) );
DFF_X1 \mreg/_11365_ ( .CK(clk ), .D(\mreg/_06504_ ), .Q(\mreg/rf[17][27] ), .QN(\mreg/_05392_ ) );
DFF_X1 \mreg/_11366_ ( .CK(clk ), .D(\mreg/_06505_ ), .Q(\mreg/rf[17][28] ), .QN(\mreg/_05391_ ) );
DFF_X1 \mreg/_11367_ ( .CK(clk ), .D(\mreg/_06506_ ), .Q(\mreg/rf[17][29] ), .QN(\mreg/_05390_ ) );
DFF_X1 \mreg/_11368_ ( .CK(clk ), .D(\mreg/_06507_ ), .Q(\mreg/rf[17][30] ), .QN(\mreg/_05389_ ) );
DFF_X1 \mreg/_11369_ ( .CK(clk ), .D(\mreg/_06508_ ), .Q(\mreg/rf[17][31] ), .QN(\mreg/_05388_ ) );
DFF_X1 \mreg/_11370_ ( .CK(clk ), .D(\mreg/_06509_ ), .Q(\mreg/rf[18][0] ), .QN(\mreg/_05387_ ) );
DFF_X1 \mreg/_11371_ ( .CK(clk ), .D(\mreg/_06510_ ), .Q(\mreg/rf[18][1] ), .QN(\mreg/_05386_ ) );
DFF_X1 \mreg/_11372_ ( .CK(clk ), .D(\mreg/_06511_ ), .Q(\mreg/rf[18][2] ), .QN(\mreg/_05385_ ) );
DFF_X1 \mreg/_11373_ ( .CK(clk ), .D(\mreg/_06512_ ), .Q(\mreg/rf[18][3] ), .QN(\mreg/_05384_ ) );
DFF_X1 \mreg/_11374_ ( .CK(clk ), .D(\mreg/_06513_ ), .Q(\mreg/rf[18][4] ), .QN(\mreg/_05383_ ) );
DFF_X1 \mreg/_11375_ ( .CK(clk ), .D(\mreg/_06514_ ), .Q(\mreg/rf[18][5] ), .QN(\mreg/_05382_ ) );
DFF_X1 \mreg/_11376_ ( .CK(clk ), .D(\mreg/_06515_ ), .Q(\mreg/rf[18][6] ), .QN(\mreg/_05381_ ) );
DFF_X1 \mreg/_11377_ ( .CK(clk ), .D(\mreg/_06516_ ), .Q(\mreg/rf[18][7] ), .QN(\mreg/_05380_ ) );
DFF_X1 \mreg/_11378_ ( .CK(clk ), .D(\mreg/_06517_ ), .Q(\mreg/rf[18][8] ), .QN(\mreg/_05379_ ) );
DFF_X1 \mreg/_11379_ ( .CK(clk ), .D(\mreg/_06518_ ), .Q(\mreg/rf[18][9] ), .QN(\mreg/_05378_ ) );
DFF_X1 \mreg/_11380_ ( .CK(clk ), .D(\mreg/_06519_ ), .Q(\mreg/rf[18][10] ), .QN(\mreg/_05377_ ) );
DFF_X1 \mreg/_11381_ ( .CK(clk ), .D(\mreg/_06520_ ), .Q(\mreg/rf[18][11] ), .QN(\mreg/_05376_ ) );
DFF_X1 \mreg/_11382_ ( .CK(clk ), .D(\mreg/_06521_ ), .Q(\mreg/rf[18][12] ), .QN(\mreg/_05375_ ) );
DFF_X1 \mreg/_11383_ ( .CK(clk ), .D(\mreg/_06522_ ), .Q(\mreg/rf[18][13] ), .QN(\mreg/_05374_ ) );
DFF_X1 \mreg/_11384_ ( .CK(clk ), .D(\mreg/_06523_ ), .Q(\mreg/rf[18][14] ), .QN(\mreg/_05373_ ) );
DFF_X1 \mreg/_11385_ ( .CK(clk ), .D(\mreg/_06524_ ), .Q(\mreg/rf[18][15] ), .QN(\mreg/_05372_ ) );
DFF_X1 \mreg/_11386_ ( .CK(clk ), .D(\mreg/_06525_ ), .Q(\mreg/rf[18][16] ), .QN(\mreg/_05371_ ) );
DFF_X1 \mreg/_11387_ ( .CK(clk ), .D(\mreg/_06526_ ), .Q(\mreg/rf[18][17] ), .QN(\mreg/_05370_ ) );
DFF_X1 \mreg/_11388_ ( .CK(clk ), .D(\mreg/_06527_ ), .Q(\mreg/rf[18][18] ), .QN(\mreg/_05369_ ) );
DFF_X1 \mreg/_11389_ ( .CK(clk ), .D(\mreg/_06528_ ), .Q(\mreg/rf[18][19] ), .QN(\mreg/_05368_ ) );
DFF_X1 \mreg/_11390_ ( .CK(clk ), .D(\mreg/_06529_ ), .Q(\mreg/rf[18][20] ), .QN(\mreg/_05367_ ) );
DFF_X1 \mreg/_11391_ ( .CK(clk ), .D(\mreg/_06530_ ), .Q(\mreg/rf[18][21] ), .QN(\mreg/_05366_ ) );
DFF_X1 \mreg/_11392_ ( .CK(clk ), .D(\mreg/_06531_ ), .Q(\mreg/rf[18][22] ), .QN(\mreg/_05365_ ) );
DFF_X1 \mreg/_11393_ ( .CK(clk ), .D(\mreg/_06532_ ), .Q(\mreg/rf[18][23] ), .QN(\mreg/_05364_ ) );
DFF_X1 \mreg/_11394_ ( .CK(clk ), .D(\mreg/_06533_ ), .Q(\mreg/rf[18][24] ), .QN(\mreg/_05363_ ) );
DFF_X1 \mreg/_11395_ ( .CK(clk ), .D(\mreg/_06534_ ), .Q(\mreg/rf[18][25] ), .QN(\mreg/_05362_ ) );
DFF_X1 \mreg/_11396_ ( .CK(clk ), .D(\mreg/_06535_ ), .Q(\mreg/rf[18][26] ), .QN(\mreg/_05361_ ) );
DFF_X1 \mreg/_11397_ ( .CK(clk ), .D(\mreg/_06536_ ), .Q(\mreg/rf[18][27] ), .QN(\mreg/_05360_ ) );
DFF_X1 \mreg/_11398_ ( .CK(clk ), .D(\mreg/_06537_ ), .Q(\mreg/rf[18][28] ), .QN(\mreg/_05359_ ) );
DFF_X1 \mreg/_11399_ ( .CK(clk ), .D(\mreg/_06538_ ), .Q(\mreg/rf[18][29] ), .QN(\mreg/_05358_ ) );
DFF_X1 \mreg/_11400_ ( .CK(clk ), .D(\mreg/_06539_ ), .Q(\mreg/rf[18][30] ), .QN(\mreg/_05357_ ) );
DFF_X1 \mreg/_11401_ ( .CK(clk ), .D(\mreg/_06540_ ), .Q(\mreg/rf[18][31] ), .QN(\mreg/_05356_ ) );
DFF_X1 \mreg/_11402_ ( .CK(clk ), .D(\mreg/_06541_ ), .Q(\mreg/rf[19][0] ), .QN(\mreg/_05355_ ) );
DFF_X1 \mreg/_11403_ ( .CK(clk ), .D(\mreg/_06542_ ), .Q(\mreg/rf[19][1] ), .QN(\mreg/_05354_ ) );
DFF_X1 \mreg/_11404_ ( .CK(clk ), .D(\mreg/_06543_ ), .Q(\mreg/rf[19][2] ), .QN(\mreg/_05353_ ) );
DFF_X1 \mreg/_11405_ ( .CK(clk ), .D(\mreg/_06544_ ), .Q(\mreg/rf[19][3] ), .QN(\mreg/_05352_ ) );
DFF_X1 \mreg/_11406_ ( .CK(clk ), .D(\mreg/_06545_ ), .Q(\mreg/rf[19][4] ), .QN(\mreg/_05351_ ) );
DFF_X1 \mreg/_11407_ ( .CK(clk ), .D(\mreg/_06546_ ), .Q(\mreg/rf[19][5] ), .QN(\mreg/_05350_ ) );
DFF_X1 \mreg/_11408_ ( .CK(clk ), .D(\mreg/_06547_ ), .Q(\mreg/rf[19][6] ), .QN(\mreg/_05349_ ) );
DFF_X1 \mreg/_11409_ ( .CK(clk ), .D(\mreg/_06548_ ), .Q(\mreg/rf[19][7] ), .QN(\mreg/_05348_ ) );
DFF_X1 \mreg/_11410_ ( .CK(clk ), .D(\mreg/_06549_ ), .Q(\mreg/rf[19][8] ), .QN(\mreg/_05347_ ) );
DFF_X1 \mreg/_11411_ ( .CK(clk ), .D(\mreg/_06550_ ), .Q(\mreg/rf[19][9] ), .QN(\mreg/_05346_ ) );
DFF_X1 \mreg/_11412_ ( .CK(clk ), .D(\mreg/_06551_ ), .Q(\mreg/rf[19][10] ), .QN(\mreg/_05345_ ) );
DFF_X1 \mreg/_11413_ ( .CK(clk ), .D(\mreg/_06552_ ), .Q(\mreg/rf[19][11] ), .QN(\mreg/_05344_ ) );
DFF_X1 \mreg/_11414_ ( .CK(clk ), .D(\mreg/_06553_ ), .Q(\mreg/rf[19][12] ), .QN(\mreg/_05343_ ) );
DFF_X1 \mreg/_11415_ ( .CK(clk ), .D(\mreg/_06554_ ), .Q(\mreg/rf[19][13] ), .QN(\mreg/_05342_ ) );
DFF_X1 \mreg/_11416_ ( .CK(clk ), .D(\mreg/_06555_ ), .Q(\mreg/rf[19][14] ), .QN(\mreg/_05341_ ) );
DFF_X1 \mreg/_11417_ ( .CK(clk ), .D(\mreg/_06556_ ), .Q(\mreg/rf[19][15] ), .QN(\mreg/_05340_ ) );
DFF_X1 \mreg/_11418_ ( .CK(clk ), .D(\mreg/_06557_ ), .Q(\mreg/rf[19][16] ), .QN(\mreg/_05339_ ) );
DFF_X1 \mreg/_11419_ ( .CK(clk ), .D(\mreg/_06558_ ), .Q(\mreg/rf[19][17] ), .QN(\mreg/_05338_ ) );
DFF_X1 \mreg/_11420_ ( .CK(clk ), .D(\mreg/_06559_ ), .Q(\mreg/rf[19][18] ), .QN(\mreg/_05337_ ) );
DFF_X1 \mreg/_11421_ ( .CK(clk ), .D(\mreg/_06560_ ), .Q(\mreg/rf[19][19] ), .QN(\mreg/_05336_ ) );
DFF_X1 \mreg/_11422_ ( .CK(clk ), .D(\mreg/_06561_ ), .Q(\mreg/rf[19][20] ), .QN(\mreg/_05335_ ) );
DFF_X1 \mreg/_11423_ ( .CK(clk ), .D(\mreg/_06562_ ), .Q(\mreg/rf[19][21] ), .QN(\mreg/_05334_ ) );
DFF_X1 \mreg/_11424_ ( .CK(clk ), .D(\mreg/_06563_ ), .Q(\mreg/rf[19][22] ), .QN(\mreg/_05333_ ) );
DFF_X1 \mreg/_11425_ ( .CK(clk ), .D(\mreg/_06564_ ), .Q(\mreg/rf[19][23] ), .QN(\mreg/_05332_ ) );
DFF_X1 \mreg/_11426_ ( .CK(clk ), .D(\mreg/_06565_ ), .Q(\mreg/rf[19][24] ), .QN(\mreg/_05331_ ) );
DFF_X1 \mreg/_11427_ ( .CK(clk ), .D(\mreg/_06566_ ), .Q(\mreg/rf[19][25] ), .QN(\mreg/_05330_ ) );
DFF_X1 \mreg/_11428_ ( .CK(clk ), .D(\mreg/_06567_ ), .Q(\mreg/rf[19][26] ), .QN(\mreg/_05329_ ) );
DFF_X1 \mreg/_11429_ ( .CK(clk ), .D(\mreg/_06568_ ), .Q(\mreg/rf[19][27] ), .QN(\mreg/_05328_ ) );
DFF_X1 \mreg/_11430_ ( .CK(clk ), .D(\mreg/_06569_ ), .Q(\mreg/rf[19][28] ), .QN(\mreg/_05327_ ) );
DFF_X1 \mreg/_11431_ ( .CK(clk ), .D(\mreg/_06570_ ), .Q(\mreg/rf[19][29] ), .QN(\mreg/_05326_ ) );
DFF_X1 \mreg/_11432_ ( .CK(clk ), .D(\mreg/_06571_ ), .Q(\mreg/rf[19][30] ), .QN(\mreg/_05325_ ) );
DFF_X1 \mreg/_11433_ ( .CK(clk ), .D(\mreg/_06572_ ), .Q(\mreg/rf[19][31] ), .QN(\mreg/_05324_ ) );
DFF_X1 \mreg/_11434_ ( .CK(clk ), .D(\mreg/_06573_ ), .Q(\mreg/rf[20][0] ), .QN(\mreg/_05323_ ) );
DFF_X1 \mreg/_11435_ ( .CK(clk ), .D(\mreg/_06574_ ), .Q(\mreg/rf[20][1] ), .QN(\mreg/_05322_ ) );
DFF_X1 \mreg/_11436_ ( .CK(clk ), .D(\mreg/_06575_ ), .Q(\mreg/rf[20][2] ), .QN(\mreg/_05321_ ) );
DFF_X1 \mreg/_11437_ ( .CK(clk ), .D(\mreg/_06576_ ), .Q(\mreg/rf[20][3] ), .QN(\mreg/_05320_ ) );
DFF_X1 \mreg/_11438_ ( .CK(clk ), .D(\mreg/_06577_ ), .Q(\mreg/rf[20][4] ), .QN(\mreg/_05319_ ) );
DFF_X1 \mreg/_11439_ ( .CK(clk ), .D(\mreg/_06578_ ), .Q(\mreg/rf[20][5] ), .QN(\mreg/_05318_ ) );
DFF_X1 \mreg/_11440_ ( .CK(clk ), .D(\mreg/_06579_ ), .Q(\mreg/rf[20][6] ), .QN(\mreg/_05317_ ) );
DFF_X1 \mreg/_11441_ ( .CK(clk ), .D(\mreg/_06580_ ), .Q(\mreg/rf[20][7] ), .QN(\mreg/_05316_ ) );
DFF_X1 \mreg/_11442_ ( .CK(clk ), .D(\mreg/_06581_ ), .Q(\mreg/rf[20][8] ), .QN(\mreg/_05315_ ) );
DFF_X1 \mreg/_11443_ ( .CK(clk ), .D(\mreg/_06582_ ), .Q(\mreg/rf[20][9] ), .QN(\mreg/_05314_ ) );
DFF_X1 \mreg/_11444_ ( .CK(clk ), .D(\mreg/_06583_ ), .Q(\mreg/rf[20][10] ), .QN(\mreg/_05313_ ) );
DFF_X1 \mreg/_11445_ ( .CK(clk ), .D(\mreg/_06584_ ), .Q(\mreg/rf[20][11] ), .QN(\mreg/_05312_ ) );
DFF_X1 \mreg/_11446_ ( .CK(clk ), .D(\mreg/_06585_ ), .Q(\mreg/rf[20][12] ), .QN(\mreg/_05311_ ) );
DFF_X1 \mreg/_11447_ ( .CK(clk ), .D(\mreg/_06586_ ), .Q(\mreg/rf[20][13] ), .QN(\mreg/_05310_ ) );
DFF_X1 \mreg/_11448_ ( .CK(clk ), .D(\mreg/_06587_ ), .Q(\mreg/rf[20][14] ), .QN(\mreg/_05309_ ) );
DFF_X1 \mreg/_11449_ ( .CK(clk ), .D(\mreg/_06588_ ), .Q(\mreg/rf[20][15] ), .QN(\mreg/_05308_ ) );
DFF_X1 \mreg/_11450_ ( .CK(clk ), .D(\mreg/_06589_ ), .Q(\mreg/rf[20][16] ), .QN(\mreg/_05307_ ) );
DFF_X1 \mreg/_11451_ ( .CK(clk ), .D(\mreg/_06590_ ), .Q(\mreg/rf[20][17] ), .QN(\mreg/_05306_ ) );
DFF_X1 \mreg/_11452_ ( .CK(clk ), .D(\mreg/_06591_ ), .Q(\mreg/rf[20][18] ), .QN(\mreg/_05305_ ) );
DFF_X1 \mreg/_11453_ ( .CK(clk ), .D(\mreg/_06592_ ), .Q(\mreg/rf[20][19] ), .QN(\mreg/_05304_ ) );
DFF_X1 \mreg/_11454_ ( .CK(clk ), .D(\mreg/_06593_ ), .Q(\mreg/rf[20][20] ), .QN(\mreg/_05303_ ) );
DFF_X1 \mreg/_11455_ ( .CK(clk ), .D(\mreg/_06594_ ), .Q(\mreg/rf[20][21] ), .QN(\mreg/_05302_ ) );
DFF_X1 \mreg/_11456_ ( .CK(clk ), .D(\mreg/_06595_ ), .Q(\mreg/rf[20][22] ), .QN(\mreg/_05301_ ) );
DFF_X1 \mreg/_11457_ ( .CK(clk ), .D(\mreg/_06596_ ), .Q(\mreg/rf[20][23] ), .QN(\mreg/_05300_ ) );
DFF_X1 \mreg/_11458_ ( .CK(clk ), .D(\mreg/_06597_ ), .Q(\mreg/rf[20][24] ), .QN(\mreg/_05299_ ) );
DFF_X1 \mreg/_11459_ ( .CK(clk ), .D(\mreg/_06598_ ), .Q(\mreg/rf[20][25] ), .QN(\mreg/_05298_ ) );
DFF_X1 \mreg/_11460_ ( .CK(clk ), .D(\mreg/_06599_ ), .Q(\mreg/rf[20][26] ), .QN(\mreg/_05297_ ) );
DFF_X1 \mreg/_11461_ ( .CK(clk ), .D(\mreg/_06600_ ), .Q(\mreg/rf[20][27] ), .QN(\mreg/_05296_ ) );
DFF_X1 \mreg/_11462_ ( .CK(clk ), .D(\mreg/_06601_ ), .Q(\mreg/rf[20][28] ), .QN(\mreg/_05295_ ) );
DFF_X1 \mreg/_11463_ ( .CK(clk ), .D(\mreg/_06602_ ), .Q(\mreg/rf[20][29] ), .QN(\mreg/_05294_ ) );
DFF_X1 \mreg/_11464_ ( .CK(clk ), .D(\mreg/_06603_ ), .Q(\mreg/rf[20][30] ), .QN(\mreg/_05293_ ) );
DFF_X1 \mreg/_11465_ ( .CK(clk ), .D(\mreg/_06604_ ), .Q(\mreg/rf[20][31] ), .QN(\mreg/_05292_ ) );
DFF_X1 \mreg/_11466_ ( .CK(clk ), .D(\mreg/_06605_ ), .Q(\mreg/rf[21][0] ), .QN(\mreg/_05291_ ) );
DFF_X1 \mreg/_11467_ ( .CK(clk ), .D(\mreg/_06606_ ), .Q(\mreg/rf[21][1] ), .QN(\mreg/_05290_ ) );
DFF_X1 \mreg/_11468_ ( .CK(clk ), .D(\mreg/_06607_ ), .Q(\mreg/rf[21][2] ), .QN(\mreg/_05289_ ) );
DFF_X1 \mreg/_11469_ ( .CK(clk ), .D(\mreg/_06608_ ), .Q(\mreg/rf[21][3] ), .QN(\mreg/_05288_ ) );
DFF_X1 \mreg/_11470_ ( .CK(clk ), .D(\mreg/_06609_ ), .Q(\mreg/rf[21][4] ), .QN(\mreg/_05287_ ) );
DFF_X1 \mreg/_11471_ ( .CK(clk ), .D(\mreg/_06610_ ), .Q(\mreg/rf[21][5] ), .QN(\mreg/_05286_ ) );
DFF_X1 \mreg/_11472_ ( .CK(clk ), .D(\mreg/_06611_ ), .Q(\mreg/rf[21][6] ), .QN(\mreg/_05285_ ) );
DFF_X1 \mreg/_11473_ ( .CK(clk ), .D(\mreg/_06612_ ), .Q(\mreg/rf[21][7] ), .QN(\mreg/_05284_ ) );
DFF_X1 \mreg/_11474_ ( .CK(clk ), .D(\mreg/_06613_ ), .Q(\mreg/rf[21][8] ), .QN(\mreg/_05283_ ) );
DFF_X1 \mreg/_11475_ ( .CK(clk ), .D(\mreg/_06614_ ), .Q(\mreg/rf[21][9] ), .QN(\mreg/_05282_ ) );
DFF_X1 \mreg/_11476_ ( .CK(clk ), .D(\mreg/_06615_ ), .Q(\mreg/rf[21][10] ), .QN(\mreg/_05281_ ) );
DFF_X1 \mreg/_11477_ ( .CK(clk ), .D(\mreg/_06616_ ), .Q(\mreg/rf[21][11] ), .QN(\mreg/_05280_ ) );
DFF_X1 \mreg/_11478_ ( .CK(clk ), .D(\mreg/_06617_ ), .Q(\mreg/rf[21][12] ), .QN(\mreg/_05279_ ) );
DFF_X1 \mreg/_11479_ ( .CK(clk ), .D(\mreg/_06618_ ), .Q(\mreg/rf[21][13] ), .QN(\mreg/_05278_ ) );
DFF_X1 \mreg/_11480_ ( .CK(clk ), .D(\mreg/_06619_ ), .Q(\mreg/rf[21][14] ), .QN(\mreg/_05277_ ) );
DFF_X1 \mreg/_11481_ ( .CK(clk ), .D(\mreg/_06620_ ), .Q(\mreg/rf[21][15] ), .QN(\mreg/_05276_ ) );
DFF_X1 \mreg/_11482_ ( .CK(clk ), .D(\mreg/_06621_ ), .Q(\mreg/rf[21][16] ), .QN(\mreg/_05275_ ) );
DFF_X1 \mreg/_11483_ ( .CK(clk ), .D(\mreg/_06622_ ), .Q(\mreg/rf[21][17] ), .QN(\mreg/_05274_ ) );
DFF_X1 \mreg/_11484_ ( .CK(clk ), .D(\mreg/_06623_ ), .Q(\mreg/rf[21][18] ), .QN(\mreg/_05273_ ) );
DFF_X1 \mreg/_11485_ ( .CK(clk ), .D(\mreg/_06624_ ), .Q(\mreg/rf[21][19] ), .QN(\mreg/_05272_ ) );
DFF_X1 \mreg/_11486_ ( .CK(clk ), .D(\mreg/_06625_ ), .Q(\mreg/rf[21][20] ), .QN(\mreg/_05271_ ) );
DFF_X1 \mreg/_11487_ ( .CK(clk ), .D(\mreg/_06626_ ), .Q(\mreg/rf[21][21] ), .QN(\mreg/_05270_ ) );
DFF_X1 \mreg/_11488_ ( .CK(clk ), .D(\mreg/_06627_ ), .Q(\mreg/rf[21][22] ), .QN(\mreg/_05269_ ) );
DFF_X1 \mreg/_11489_ ( .CK(clk ), .D(\mreg/_06628_ ), .Q(\mreg/rf[21][23] ), .QN(\mreg/_05268_ ) );
DFF_X1 \mreg/_11490_ ( .CK(clk ), .D(\mreg/_06629_ ), .Q(\mreg/rf[21][24] ), .QN(\mreg/_05267_ ) );
DFF_X1 \mreg/_11491_ ( .CK(clk ), .D(\mreg/_06630_ ), .Q(\mreg/rf[21][25] ), .QN(\mreg/_05266_ ) );
DFF_X1 \mreg/_11492_ ( .CK(clk ), .D(\mreg/_06631_ ), .Q(\mreg/rf[21][26] ), .QN(\mreg/_05265_ ) );
DFF_X1 \mreg/_11493_ ( .CK(clk ), .D(\mreg/_06632_ ), .Q(\mreg/rf[21][27] ), .QN(\mreg/_05264_ ) );
DFF_X1 \mreg/_11494_ ( .CK(clk ), .D(\mreg/_06633_ ), .Q(\mreg/rf[21][28] ), .QN(\mreg/_05263_ ) );
DFF_X1 \mreg/_11495_ ( .CK(clk ), .D(\mreg/_06634_ ), .Q(\mreg/rf[21][29] ), .QN(\mreg/_05262_ ) );
DFF_X1 \mreg/_11496_ ( .CK(clk ), .D(\mreg/_06635_ ), .Q(\mreg/rf[21][30] ), .QN(\mreg/_05261_ ) );
DFF_X1 \mreg/_11497_ ( .CK(clk ), .D(\mreg/_06636_ ), .Q(\mreg/rf[21][31] ), .QN(\mreg/_05260_ ) );
DFF_X1 \mreg/_11498_ ( .CK(clk ), .D(\mreg/_06637_ ), .Q(\mreg/rf[22][0] ), .QN(\mreg/_05259_ ) );
DFF_X1 \mreg/_11499_ ( .CK(clk ), .D(\mreg/_06638_ ), .Q(\mreg/rf[22][1] ), .QN(\mreg/_05258_ ) );
DFF_X1 \mreg/_11500_ ( .CK(clk ), .D(\mreg/_06639_ ), .Q(\mreg/rf[22][2] ), .QN(\mreg/_05257_ ) );
DFF_X1 \mreg/_11501_ ( .CK(clk ), .D(\mreg/_06640_ ), .Q(\mreg/rf[22][3] ), .QN(\mreg/_05256_ ) );
DFF_X1 \mreg/_11502_ ( .CK(clk ), .D(\mreg/_06641_ ), .Q(\mreg/rf[22][4] ), .QN(\mreg/_05255_ ) );
DFF_X1 \mreg/_11503_ ( .CK(clk ), .D(\mreg/_06642_ ), .Q(\mreg/rf[22][5] ), .QN(\mreg/_05254_ ) );
DFF_X1 \mreg/_11504_ ( .CK(clk ), .D(\mreg/_06643_ ), .Q(\mreg/rf[22][6] ), .QN(\mreg/_05253_ ) );
DFF_X1 \mreg/_11505_ ( .CK(clk ), .D(\mreg/_06644_ ), .Q(\mreg/rf[22][7] ), .QN(\mreg/_05252_ ) );
DFF_X1 \mreg/_11506_ ( .CK(clk ), .D(\mreg/_06645_ ), .Q(\mreg/rf[22][8] ), .QN(\mreg/_05251_ ) );
DFF_X1 \mreg/_11507_ ( .CK(clk ), .D(\mreg/_06646_ ), .Q(\mreg/rf[22][9] ), .QN(\mreg/_05250_ ) );
DFF_X1 \mreg/_11508_ ( .CK(clk ), .D(\mreg/_06647_ ), .Q(\mreg/rf[22][10] ), .QN(\mreg/_05249_ ) );
DFF_X1 \mreg/_11509_ ( .CK(clk ), .D(\mreg/_06648_ ), .Q(\mreg/rf[22][11] ), .QN(\mreg/_05248_ ) );
DFF_X1 \mreg/_11510_ ( .CK(clk ), .D(\mreg/_06649_ ), .Q(\mreg/rf[22][12] ), .QN(\mreg/_05247_ ) );
DFF_X1 \mreg/_11511_ ( .CK(clk ), .D(\mreg/_06650_ ), .Q(\mreg/rf[22][13] ), .QN(\mreg/_05246_ ) );
DFF_X1 \mreg/_11512_ ( .CK(clk ), .D(\mreg/_06651_ ), .Q(\mreg/rf[22][14] ), .QN(\mreg/_05245_ ) );
DFF_X1 \mreg/_11513_ ( .CK(clk ), .D(\mreg/_06652_ ), .Q(\mreg/rf[22][15] ), .QN(\mreg/_05244_ ) );
DFF_X1 \mreg/_11514_ ( .CK(clk ), .D(\mreg/_06653_ ), .Q(\mreg/rf[22][16] ), .QN(\mreg/_05243_ ) );
DFF_X1 \mreg/_11515_ ( .CK(clk ), .D(\mreg/_06654_ ), .Q(\mreg/rf[22][17] ), .QN(\mreg/_05242_ ) );
DFF_X1 \mreg/_11516_ ( .CK(clk ), .D(\mreg/_06655_ ), .Q(\mreg/rf[22][18] ), .QN(\mreg/_05241_ ) );
DFF_X1 \mreg/_11517_ ( .CK(clk ), .D(\mreg/_06656_ ), .Q(\mreg/rf[22][19] ), .QN(\mreg/_05240_ ) );
DFF_X1 \mreg/_11518_ ( .CK(clk ), .D(\mreg/_06657_ ), .Q(\mreg/rf[22][20] ), .QN(\mreg/_05239_ ) );
DFF_X1 \mreg/_11519_ ( .CK(clk ), .D(\mreg/_06658_ ), .Q(\mreg/rf[22][21] ), .QN(\mreg/_05238_ ) );
DFF_X1 \mreg/_11520_ ( .CK(clk ), .D(\mreg/_06659_ ), .Q(\mreg/rf[22][22] ), .QN(\mreg/_05237_ ) );
DFF_X1 \mreg/_11521_ ( .CK(clk ), .D(\mreg/_06660_ ), .Q(\mreg/rf[22][23] ), .QN(\mreg/_05236_ ) );
DFF_X1 \mreg/_11522_ ( .CK(clk ), .D(\mreg/_06661_ ), .Q(\mreg/rf[22][24] ), .QN(\mreg/_05235_ ) );
DFF_X1 \mreg/_11523_ ( .CK(clk ), .D(\mreg/_06662_ ), .Q(\mreg/rf[22][25] ), .QN(\mreg/_05234_ ) );
DFF_X1 \mreg/_11524_ ( .CK(clk ), .D(\mreg/_06663_ ), .Q(\mreg/rf[22][26] ), .QN(\mreg/_05233_ ) );
DFF_X1 \mreg/_11525_ ( .CK(clk ), .D(\mreg/_06664_ ), .Q(\mreg/rf[22][27] ), .QN(\mreg/_05232_ ) );
DFF_X1 \mreg/_11526_ ( .CK(clk ), .D(\mreg/_06665_ ), .Q(\mreg/rf[22][28] ), .QN(\mreg/_05231_ ) );
DFF_X1 \mreg/_11527_ ( .CK(clk ), .D(\mreg/_06666_ ), .Q(\mreg/rf[22][29] ), .QN(\mreg/_05230_ ) );
DFF_X1 \mreg/_11528_ ( .CK(clk ), .D(\mreg/_06667_ ), .Q(\mreg/rf[22][30] ), .QN(\mreg/_05229_ ) );
DFF_X1 \mreg/_11529_ ( .CK(clk ), .D(\mreg/_06668_ ), .Q(\mreg/rf[22][31] ), .QN(\mreg/_05228_ ) );
DFF_X1 \mreg/_11530_ ( .CK(clk ), .D(\mreg/_06669_ ), .Q(\mreg/rf[23][0] ), .QN(\mreg/_05227_ ) );
DFF_X1 \mreg/_11531_ ( .CK(clk ), .D(\mreg/_06670_ ), .Q(\mreg/rf[23][1] ), .QN(\mreg/_05226_ ) );
DFF_X1 \mreg/_11532_ ( .CK(clk ), .D(\mreg/_06671_ ), .Q(\mreg/rf[23][2] ), .QN(\mreg/_05225_ ) );
DFF_X1 \mreg/_11533_ ( .CK(clk ), .D(\mreg/_06672_ ), .Q(\mreg/rf[23][3] ), .QN(\mreg/_05224_ ) );
DFF_X1 \mreg/_11534_ ( .CK(clk ), .D(\mreg/_06673_ ), .Q(\mreg/rf[23][4] ), .QN(\mreg/_05223_ ) );
DFF_X1 \mreg/_11535_ ( .CK(clk ), .D(\mreg/_06674_ ), .Q(\mreg/rf[23][5] ), .QN(\mreg/_05222_ ) );
DFF_X1 \mreg/_11536_ ( .CK(clk ), .D(\mreg/_06675_ ), .Q(\mreg/rf[23][6] ), .QN(\mreg/_05221_ ) );
DFF_X1 \mreg/_11537_ ( .CK(clk ), .D(\mreg/_06676_ ), .Q(\mreg/rf[23][7] ), .QN(\mreg/_05220_ ) );
DFF_X1 \mreg/_11538_ ( .CK(clk ), .D(\mreg/_06677_ ), .Q(\mreg/rf[23][8] ), .QN(\mreg/_05219_ ) );
DFF_X1 \mreg/_11539_ ( .CK(clk ), .D(\mreg/_06678_ ), .Q(\mreg/rf[23][9] ), .QN(\mreg/_05218_ ) );
DFF_X1 \mreg/_11540_ ( .CK(clk ), .D(\mreg/_06679_ ), .Q(\mreg/rf[23][10] ), .QN(\mreg/_05217_ ) );
DFF_X1 \mreg/_11541_ ( .CK(clk ), .D(\mreg/_06680_ ), .Q(\mreg/rf[23][11] ), .QN(\mreg/_05216_ ) );
DFF_X1 \mreg/_11542_ ( .CK(clk ), .D(\mreg/_06681_ ), .Q(\mreg/rf[23][12] ), .QN(\mreg/_05215_ ) );
DFF_X1 \mreg/_11543_ ( .CK(clk ), .D(\mreg/_06682_ ), .Q(\mreg/rf[23][13] ), .QN(\mreg/_05214_ ) );
DFF_X1 \mreg/_11544_ ( .CK(clk ), .D(\mreg/_06683_ ), .Q(\mreg/rf[23][14] ), .QN(\mreg/_05213_ ) );
DFF_X1 \mreg/_11545_ ( .CK(clk ), .D(\mreg/_06684_ ), .Q(\mreg/rf[23][15] ), .QN(\mreg/_05212_ ) );
DFF_X1 \mreg/_11546_ ( .CK(clk ), .D(\mreg/_06685_ ), .Q(\mreg/rf[23][16] ), .QN(\mreg/_05211_ ) );
DFF_X1 \mreg/_11547_ ( .CK(clk ), .D(\mreg/_06686_ ), .Q(\mreg/rf[23][17] ), .QN(\mreg/_05210_ ) );
DFF_X1 \mreg/_11548_ ( .CK(clk ), .D(\mreg/_06687_ ), .Q(\mreg/rf[23][18] ), .QN(\mreg/_05209_ ) );
DFF_X1 \mreg/_11549_ ( .CK(clk ), .D(\mreg/_06688_ ), .Q(\mreg/rf[23][19] ), .QN(\mreg/_05208_ ) );
DFF_X1 \mreg/_11550_ ( .CK(clk ), .D(\mreg/_06689_ ), .Q(\mreg/rf[23][20] ), .QN(\mreg/_05207_ ) );
DFF_X1 \mreg/_11551_ ( .CK(clk ), .D(\mreg/_06690_ ), .Q(\mreg/rf[23][21] ), .QN(\mreg/_05206_ ) );
DFF_X1 \mreg/_11552_ ( .CK(clk ), .D(\mreg/_06691_ ), .Q(\mreg/rf[23][22] ), .QN(\mreg/_05205_ ) );
DFF_X1 \mreg/_11553_ ( .CK(clk ), .D(\mreg/_06692_ ), .Q(\mreg/rf[23][23] ), .QN(\mreg/_05204_ ) );
DFF_X1 \mreg/_11554_ ( .CK(clk ), .D(\mreg/_06693_ ), .Q(\mreg/rf[23][24] ), .QN(\mreg/_05203_ ) );
DFF_X1 \mreg/_11555_ ( .CK(clk ), .D(\mreg/_06694_ ), .Q(\mreg/rf[23][25] ), .QN(\mreg/_05202_ ) );
DFF_X1 \mreg/_11556_ ( .CK(clk ), .D(\mreg/_06695_ ), .Q(\mreg/rf[23][26] ), .QN(\mreg/_05201_ ) );
DFF_X1 \mreg/_11557_ ( .CK(clk ), .D(\mreg/_06696_ ), .Q(\mreg/rf[23][27] ), .QN(\mreg/_05200_ ) );
DFF_X1 \mreg/_11558_ ( .CK(clk ), .D(\mreg/_06697_ ), .Q(\mreg/rf[23][28] ), .QN(\mreg/_05199_ ) );
DFF_X1 \mreg/_11559_ ( .CK(clk ), .D(\mreg/_06698_ ), .Q(\mreg/rf[23][29] ), .QN(\mreg/_05198_ ) );
DFF_X1 \mreg/_11560_ ( .CK(clk ), .D(\mreg/_06699_ ), .Q(\mreg/rf[23][30] ), .QN(\mreg/_05197_ ) );
DFF_X1 \mreg/_11561_ ( .CK(clk ), .D(\mreg/_06700_ ), .Q(\mreg/rf[23][31] ), .QN(\mreg/_05196_ ) );
DFF_X1 \mreg/_11562_ ( .CK(clk ), .D(\mreg/_06701_ ), .Q(\mreg/rf[24][0] ), .QN(\mreg/_05195_ ) );
DFF_X1 \mreg/_11563_ ( .CK(clk ), .D(\mreg/_06702_ ), .Q(\mreg/rf[24][1] ), .QN(\mreg/_05194_ ) );
DFF_X1 \mreg/_11564_ ( .CK(clk ), .D(\mreg/_06703_ ), .Q(\mreg/rf[24][2] ), .QN(\mreg/_05193_ ) );
DFF_X1 \mreg/_11565_ ( .CK(clk ), .D(\mreg/_06704_ ), .Q(\mreg/rf[24][3] ), .QN(\mreg/_05192_ ) );
DFF_X1 \mreg/_11566_ ( .CK(clk ), .D(\mreg/_06705_ ), .Q(\mreg/rf[24][4] ), .QN(\mreg/_05191_ ) );
DFF_X1 \mreg/_11567_ ( .CK(clk ), .D(\mreg/_06706_ ), .Q(\mreg/rf[24][5] ), .QN(\mreg/_05190_ ) );
DFF_X1 \mreg/_11568_ ( .CK(clk ), .D(\mreg/_06707_ ), .Q(\mreg/rf[24][6] ), .QN(\mreg/_05189_ ) );
DFF_X1 \mreg/_11569_ ( .CK(clk ), .D(\mreg/_06708_ ), .Q(\mreg/rf[24][7] ), .QN(\mreg/_05188_ ) );
DFF_X1 \mreg/_11570_ ( .CK(clk ), .D(\mreg/_06709_ ), .Q(\mreg/rf[24][8] ), .QN(\mreg/_05187_ ) );
DFF_X1 \mreg/_11571_ ( .CK(clk ), .D(\mreg/_06710_ ), .Q(\mreg/rf[24][9] ), .QN(\mreg/_05186_ ) );
DFF_X1 \mreg/_11572_ ( .CK(clk ), .D(\mreg/_06711_ ), .Q(\mreg/rf[24][10] ), .QN(\mreg/_05185_ ) );
DFF_X1 \mreg/_11573_ ( .CK(clk ), .D(\mreg/_06712_ ), .Q(\mreg/rf[24][11] ), .QN(\mreg/_05184_ ) );
DFF_X1 \mreg/_11574_ ( .CK(clk ), .D(\mreg/_06713_ ), .Q(\mreg/rf[24][12] ), .QN(\mreg/_05183_ ) );
DFF_X1 \mreg/_11575_ ( .CK(clk ), .D(\mreg/_06714_ ), .Q(\mreg/rf[24][13] ), .QN(\mreg/_05182_ ) );
DFF_X1 \mreg/_11576_ ( .CK(clk ), .D(\mreg/_06715_ ), .Q(\mreg/rf[24][14] ), .QN(\mreg/_05181_ ) );
DFF_X1 \mreg/_11577_ ( .CK(clk ), .D(\mreg/_06716_ ), .Q(\mreg/rf[24][15] ), .QN(\mreg/_05180_ ) );
DFF_X1 \mreg/_11578_ ( .CK(clk ), .D(\mreg/_06717_ ), .Q(\mreg/rf[24][16] ), .QN(\mreg/_05179_ ) );
DFF_X1 \mreg/_11579_ ( .CK(clk ), .D(\mreg/_06718_ ), .Q(\mreg/rf[24][17] ), .QN(\mreg/_05178_ ) );
DFF_X1 \mreg/_11580_ ( .CK(clk ), .D(\mreg/_06719_ ), .Q(\mreg/rf[24][18] ), .QN(\mreg/_05177_ ) );
DFF_X1 \mreg/_11581_ ( .CK(clk ), .D(\mreg/_06720_ ), .Q(\mreg/rf[24][19] ), .QN(\mreg/_05176_ ) );
DFF_X1 \mreg/_11582_ ( .CK(clk ), .D(\mreg/_06721_ ), .Q(\mreg/rf[24][20] ), .QN(\mreg/_05175_ ) );
DFF_X1 \mreg/_11583_ ( .CK(clk ), .D(\mreg/_06722_ ), .Q(\mreg/rf[24][21] ), .QN(\mreg/_05174_ ) );
DFF_X1 \mreg/_11584_ ( .CK(clk ), .D(\mreg/_06723_ ), .Q(\mreg/rf[24][22] ), .QN(\mreg/_05173_ ) );
DFF_X1 \mreg/_11585_ ( .CK(clk ), .D(\mreg/_06724_ ), .Q(\mreg/rf[24][23] ), .QN(\mreg/_05172_ ) );
DFF_X1 \mreg/_11586_ ( .CK(clk ), .D(\mreg/_06725_ ), .Q(\mreg/rf[24][24] ), .QN(\mreg/_05171_ ) );
DFF_X1 \mreg/_11587_ ( .CK(clk ), .D(\mreg/_06726_ ), .Q(\mreg/rf[24][25] ), .QN(\mreg/_05170_ ) );
DFF_X1 \mreg/_11588_ ( .CK(clk ), .D(\mreg/_06727_ ), .Q(\mreg/rf[24][26] ), .QN(\mreg/_05169_ ) );
DFF_X1 \mreg/_11589_ ( .CK(clk ), .D(\mreg/_06728_ ), .Q(\mreg/rf[24][27] ), .QN(\mreg/_05168_ ) );
DFF_X1 \mreg/_11590_ ( .CK(clk ), .D(\mreg/_06729_ ), .Q(\mreg/rf[24][28] ), .QN(\mreg/_05167_ ) );
DFF_X1 \mreg/_11591_ ( .CK(clk ), .D(\mreg/_06730_ ), .Q(\mreg/rf[24][29] ), .QN(\mreg/_05166_ ) );
DFF_X1 \mreg/_11592_ ( .CK(clk ), .D(\mreg/_06731_ ), .Q(\mreg/rf[24][30] ), .QN(\mreg/_05165_ ) );
DFF_X1 \mreg/_11593_ ( .CK(clk ), .D(\mreg/_06732_ ), .Q(\mreg/rf[24][31] ), .QN(\mreg/_05164_ ) );
DFF_X1 \mreg/_11594_ ( .CK(clk ), .D(\mreg/_06733_ ), .Q(\mreg/rf[25][0] ), .QN(\mreg/_05163_ ) );
DFF_X1 \mreg/_11595_ ( .CK(clk ), .D(\mreg/_06734_ ), .Q(\mreg/rf[25][1] ), .QN(\mreg/_05162_ ) );
DFF_X1 \mreg/_11596_ ( .CK(clk ), .D(\mreg/_06735_ ), .Q(\mreg/rf[25][2] ), .QN(\mreg/_05161_ ) );
DFF_X1 \mreg/_11597_ ( .CK(clk ), .D(\mreg/_06736_ ), .Q(\mreg/rf[25][3] ), .QN(\mreg/_05160_ ) );
DFF_X1 \mreg/_11598_ ( .CK(clk ), .D(\mreg/_06737_ ), .Q(\mreg/rf[25][4] ), .QN(\mreg/_05159_ ) );
DFF_X1 \mreg/_11599_ ( .CK(clk ), .D(\mreg/_06738_ ), .Q(\mreg/rf[25][5] ), .QN(\mreg/_05158_ ) );
DFF_X1 \mreg/_11600_ ( .CK(clk ), .D(\mreg/_06739_ ), .Q(\mreg/rf[25][6] ), .QN(\mreg/_05157_ ) );
DFF_X1 \mreg/_11601_ ( .CK(clk ), .D(\mreg/_06740_ ), .Q(\mreg/rf[25][7] ), .QN(\mreg/_05156_ ) );
DFF_X1 \mreg/_11602_ ( .CK(clk ), .D(\mreg/_06741_ ), .Q(\mreg/rf[25][8] ), .QN(\mreg/_05155_ ) );
DFF_X1 \mreg/_11603_ ( .CK(clk ), .D(\mreg/_06742_ ), .Q(\mreg/rf[25][9] ), .QN(\mreg/_05154_ ) );
DFF_X1 \mreg/_11604_ ( .CK(clk ), .D(\mreg/_06743_ ), .Q(\mreg/rf[25][10] ), .QN(\mreg/_05153_ ) );
DFF_X1 \mreg/_11605_ ( .CK(clk ), .D(\mreg/_06744_ ), .Q(\mreg/rf[25][11] ), .QN(\mreg/_05152_ ) );
DFF_X1 \mreg/_11606_ ( .CK(clk ), .D(\mreg/_06745_ ), .Q(\mreg/rf[25][12] ), .QN(\mreg/_05151_ ) );
DFF_X1 \mreg/_11607_ ( .CK(clk ), .D(\mreg/_06746_ ), .Q(\mreg/rf[25][13] ), .QN(\mreg/_05150_ ) );
DFF_X1 \mreg/_11608_ ( .CK(clk ), .D(\mreg/_06747_ ), .Q(\mreg/rf[25][14] ), .QN(\mreg/_05149_ ) );
DFF_X1 \mreg/_11609_ ( .CK(clk ), .D(\mreg/_06748_ ), .Q(\mreg/rf[25][15] ), .QN(\mreg/_05148_ ) );
DFF_X1 \mreg/_11610_ ( .CK(clk ), .D(\mreg/_06749_ ), .Q(\mreg/rf[25][16] ), .QN(\mreg/_05147_ ) );
DFF_X1 \mreg/_11611_ ( .CK(clk ), .D(\mreg/_06750_ ), .Q(\mreg/rf[25][17] ), .QN(\mreg/_05146_ ) );
DFF_X1 \mreg/_11612_ ( .CK(clk ), .D(\mreg/_06751_ ), .Q(\mreg/rf[25][18] ), .QN(\mreg/_05145_ ) );
DFF_X1 \mreg/_11613_ ( .CK(clk ), .D(\mreg/_06752_ ), .Q(\mreg/rf[25][19] ), .QN(\mreg/_05144_ ) );
DFF_X1 \mreg/_11614_ ( .CK(clk ), .D(\mreg/_06753_ ), .Q(\mreg/rf[25][20] ), .QN(\mreg/_05143_ ) );
DFF_X1 \mreg/_11615_ ( .CK(clk ), .D(\mreg/_06754_ ), .Q(\mreg/rf[25][21] ), .QN(\mreg/_05142_ ) );
DFF_X1 \mreg/_11616_ ( .CK(clk ), .D(\mreg/_06755_ ), .Q(\mreg/rf[25][22] ), .QN(\mreg/_05141_ ) );
DFF_X1 \mreg/_11617_ ( .CK(clk ), .D(\mreg/_06756_ ), .Q(\mreg/rf[25][23] ), .QN(\mreg/_05140_ ) );
DFF_X1 \mreg/_11618_ ( .CK(clk ), .D(\mreg/_06757_ ), .Q(\mreg/rf[25][24] ), .QN(\mreg/_05139_ ) );
DFF_X1 \mreg/_11619_ ( .CK(clk ), .D(\mreg/_06758_ ), .Q(\mreg/rf[25][25] ), .QN(\mreg/_05138_ ) );
DFF_X1 \mreg/_11620_ ( .CK(clk ), .D(\mreg/_06759_ ), .Q(\mreg/rf[25][26] ), .QN(\mreg/_05137_ ) );
DFF_X1 \mreg/_11621_ ( .CK(clk ), .D(\mreg/_06760_ ), .Q(\mreg/rf[25][27] ), .QN(\mreg/_05136_ ) );
DFF_X1 \mreg/_11622_ ( .CK(clk ), .D(\mreg/_06761_ ), .Q(\mreg/rf[25][28] ), .QN(\mreg/_05135_ ) );
DFF_X1 \mreg/_11623_ ( .CK(clk ), .D(\mreg/_06762_ ), .Q(\mreg/rf[25][29] ), .QN(\mreg/_05134_ ) );
DFF_X1 \mreg/_11624_ ( .CK(clk ), .D(\mreg/_06763_ ), .Q(\mreg/rf[25][30] ), .QN(\mreg/_05133_ ) );
DFF_X1 \mreg/_11625_ ( .CK(clk ), .D(\mreg/_06764_ ), .Q(\mreg/rf[25][31] ), .QN(\mreg/_05132_ ) );
DFF_X1 \mreg/_11626_ ( .CK(clk ), .D(\mreg/_06765_ ), .Q(\mreg/rf[26][0] ), .QN(\mreg/_05131_ ) );
DFF_X1 \mreg/_11627_ ( .CK(clk ), .D(\mreg/_06766_ ), .Q(\mreg/rf[26][1] ), .QN(\mreg/_05130_ ) );
DFF_X1 \mreg/_11628_ ( .CK(clk ), .D(\mreg/_06767_ ), .Q(\mreg/rf[26][2] ), .QN(\mreg/_05129_ ) );
DFF_X1 \mreg/_11629_ ( .CK(clk ), .D(\mreg/_06768_ ), .Q(\mreg/rf[26][3] ), .QN(\mreg/_05128_ ) );
DFF_X1 \mreg/_11630_ ( .CK(clk ), .D(\mreg/_06769_ ), .Q(\mreg/rf[26][4] ), .QN(\mreg/_05127_ ) );
DFF_X1 \mreg/_11631_ ( .CK(clk ), .D(\mreg/_06770_ ), .Q(\mreg/rf[26][5] ), .QN(\mreg/_05126_ ) );
DFF_X1 \mreg/_11632_ ( .CK(clk ), .D(\mreg/_06771_ ), .Q(\mreg/rf[26][6] ), .QN(\mreg/_05125_ ) );
DFF_X1 \mreg/_11633_ ( .CK(clk ), .D(\mreg/_06772_ ), .Q(\mreg/rf[26][7] ), .QN(\mreg/_05124_ ) );
DFF_X1 \mreg/_11634_ ( .CK(clk ), .D(\mreg/_06773_ ), .Q(\mreg/rf[26][8] ), .QN(\mreg/_05123_ ) );
DFF_X1 \mreg/_11635_ ( .CK(clk ), .D(\mreg/_06774_ ), .Q(\mreg/rf[26][9] ), .QN(\mreg/_05122_ ) );
DFF_X1 \mreg/_11636_ ( .CK(clk ), .D(\mreg/_06775_ ), .Q(\mreg/rf[26][10] ), .QN(\mreg/_05121_ ) );
DFF_X1 \mreg/_11637_ ( .CK(clk ), .D(\mreg/_06776_ ), .Q(\mreg/rf[26][11] ), .QN(\mreg/_05120_ ) );
DFF_X1 \mreg/_11638_ ( .CK(clk ), .D(\mreg/_06777_ ), .Q(\mreg/rf[26][12] ), .QN(\mreg/_05119_ ) );
DFF_X1 \mreg/_11639_ ( .CK(clk ), .D(\mreg/_06778_ ), .Q(\mreg/rf[26][13] ), .QN(\mreg/_05118_ ) );
DFF_X1 \mreg/_11640_ ( .CK(clk ), .D(\mreg/_06779_ ), .Q(\mreg/rf[26][14] ), .QN(\mreg/_05117_ ) );
DFF_X1 \mreg/_11641_ ( .CK(clk ), .D(\mreg/_06780_ ), .Q(\mreg/rf[26][15] ), .QN(\mreg/_05116_ ) );
DFF_X1 \mreg/_11642_ ( .CK(clk ), .D(\mreg/_06781_ ), .Q(\mreg/rf[26][16] ), .QN(\mreg/_05115_ ) );
DFF_X1 \mreg/_11643_ ( .CK(clk ), .D(\mreg/_06782_ ), .Q(\mreg/rf[26][17] ), .QN(\mreg/_05114_ ) );
DFF_X1 \mreg/_11644_ ( .CK(clk ), .D(\mreg/_06783_ ), .Q(\mreg/rf[26][18] ), .QN(\mreg/_05113_ ) );
DFF_X1 \mreg/_11645_ ( .CK(clk ), .D(\mreg/_06784_ ), .Q(\mreg/rf[26][19] ), .QN(\mreg/_05112_ ) );
DFF_X1 \mreg/_11646_ ( .CK(clk ), .D(\mreg/_06785_ ), .Q(\mreg/rf[26][20] ), .QN(\mreg/_05111_ ) );
DFF_X1 \mreg/_11647_ ( .CK(clk ), .D(\mreg/_06786_ ), .Q(\mreg/rf[26][21] ), .QN(\mreg/_05110_ ) );
DFF_X1 \mreg/_11648_ ( .CK(clk ), .D(\mreg/_06787_ ), .Q(\mreg/rf[26][22] ), .QN(\mreg/_05109_ ) );
DFF_X1 \mreg/_11649_ ( .CK(clk ), .D(\mreg/_06788_ ), .Q(\mreg/rf[26][23] ), .QN(\mreg/_05108_ ) );
DFF_X1 \mreg/_11650_ ( .CK(clk ), .D(\mreg/_06789_ ), .Q(\mreg/rf[26][24] ), .QN(\mreg/_05107_ ) );
DFF_X1 \mreg/_11651_ ( .CK(clk ), .D(\mreg/_06790_ ), .Q(\mreg/rf[26][25] ), .QN(\mreg/_05106_ ) );
DFF_X1 \mreg/_11652_ ( .CK(clk ), .D(\mreg/_06791_ ), .Q(\mreg/rf[26][26] ), .QN(\mreg/_05105_ ) );
DFF_X1 \mreg/_11653_ ( .CK(clk ), .D(\mreg/_06792_ ), .Q(\mreg/rf[26][27] ), .QN(\mreg/_05104_ ) );
DFF_X1 \mreg/_11654_ ( .CK(clk ), .D(\mreg/_06793_ ), .Q(\mreg/rf[26][28] ), .QN(\mreg/_05103_ ) );
DFF_X1 \mreg/_11655_ ( .CK(clk ), .D(\mreg/_06794_ ), .Q(\mreg/rf[26][29] ), .QN(\mreg/_05102_ ) );
DFF_X1 \mreg/_11656_ ( .CK(clk ), .D(\mreg/_06795_ ), .Q(\mreg/rf[26][30] ), .QN(\mreg/_05101_ ) );
DFF_X1 \mreg/_11657_ ( .CK(clk ), .D(\mreg/_06796_ ), .Q(\mreg/rf[26][31] ), .QN(\mreg/_05100_ ) );
DFF_X1 \mreg/_11658_ ( .CK(clk ), .D(\mreg/_06797_ ), .Q(\mreg/rf[27][0] ), .QN(\mreg/_05099_ ) );
DFF_X1 \mreg/_11659_ ( .CK(clk ), .D(\mreg/_06798_ ), .Q(\mreg/rf[27][1] ), .QN(\mreg/_05098_ ) );
DFF_X1 \mreg/_11660_ ( .CK(clk ), .D(\mreg/_06799_ ), .Q(\mreg/rf[27][2] ), .QN(\mreg/_05097_ ) );
DFF_X1 \mreg/_11661_ ( .CK(clk ), .D(\mreg/_06800_ ), .Q(\mreg/rf[27][3] ), .QN(\mreg/_05096_ ) );
DFF_X1 \mreg/_11662_ ( .CK(clk ), .D(\mreg/_06801_ ), .Q(\mreg/rf[27][4] ), .QN(\mreg/_05095_ ) );
DFF_X1 \mreg/_11663_ ( .CK(clk ), .D(\mreg/_06802_ ), .Q(\mreg/rf[27][5] ), .QN(\mreg/_05094_ ) );
DFF_X1 \mreg/_11664_ ( .CK(clk ), .D(\mreg/_06803_ ), .Q(\mreg/rf[27][6] ), .QN(\mreg/_05093_ ) );
DFF_X1 \mreg/_11665_ ( .CK(clk ), .D(\mreg/_06804_ ), .Q(\mreg/rf[27][7] ), .QN(\mreg/_05092_ ) );
DFF_X1 \mreg/_11666_ ( .CK(clk ), .D(\mreg/_06805_ ), .Q(\mreg/rf[27][8] ), .QN(\mreg/_05091_ ) );
DFF_X1 \mreg/_11667_ ( .CK(clk ), .D(\mreg/_06806_ ), .Q(\mreg/rf[27][9] ), .QN(\mreg/_05090_ ) );
DFF_X1 \mreg/_11668_ ( .CK(clk ), .D(\mreg/_06807_ ), .Q(\mreg/rf[27][10] ), .QN(\mreg/_05089_ ) );
DFF_X1 \mreg/_11669_ ( .CK(clk ), .D(\mreg/_06808_ ), .Q(\mreg/rf[27][11] ), .QN(\mreg/_05088_ ) );
DFF_X1 \mreg/_11670_ ( .CK(clk ), .D(\mreg/_06809_ ), .Q(\mreg/rf[27][12] ), .QN(\mreg/_05087_ ) );
DFF_X1 \mreg/_11671_ ( .CK(clk ), .D(\mreg/_06810_ ), .Q(\mreg/rf[27][13] ), .QN(\mreg/_05086_ ) );
DFF_X1 \mreg/_11672_ ( .CK(clk ), .D(\mreg/_06811_ ), .Q(\mreg/rf[27][14] ), .QN(\mreg/_05085_ ) );
DFF_X1 \mreg/_11673_ ( .CK(clk ), .D(\mreg/_06812_ ), .Q(\mreg/rf[27][15] ), .QN(\mreg/_05084_ ) );
DFF_X1 \mreg/_11674_ ( .CK(clk ), .D(\mreg/_06813_ ), .Q(\mreg/rf[27][16] ), .QN(\mreg/_05083_ ) );
DFF_X1 \mreg/_11675_ ( .CK(clk ), .D(\mreg/_06814_ ), .Q(\mreg/rf[27][17] ), .QN(\mreg/_05082_ ) );
DFF_X1 \mreg/_11676_ ( .CK(clk ), .D(\mreg/_06815_ ), .Q(\mreg/rf[27][18] ), .QN(\mreg/_05081_ ) );
DFF_X1 \mreg/_11677_ ( .CK(clk ), .D(\mreg/_06816_ ), .Q(\mreg/rf[27][19] ), .QN(\mreg/_05080_ ) );
DFF_X1 \mreg/_11678_ ( .CK(clk ), .D(\mreg/_06817_ ), .Q(\mreg/rf[27][20] ), .QN(\mreg/_05079_ ) );
DFF_X1 \mreg/_11679_ ( .CK(clk ), .D(\mreg/_06818_ ), .Q(\mreg/rf[27][21] ), .QN(\mreg/_05078_ ) );
DFF_X1 \mreg/_11680_ ( .CK(clk ), .D(\mreg/_06819_ ), .Q(\mreg/rf[27][22] ), .QN(\mreg/_05077_ ) );
DFF_X1 \mreg/_11681_ ( .CK(clk ), .D(\mreg/_06820_ ), .Q(\mreg/rf[27][23] ), .QN(\mreg/_05076_ ) );
DFF_X1 \mreg/_11682_ ( .CK(clk ), .D(\mreg/_06821_ ), .Q(\mreg/rf[27][24] ), .QN(\mreg/_05075_ ) );
DFF_X1 \mreg/_11683_ ( .CK(clk ), .D(\mreg/_06822_ ), .Q(\mreg/rf[27][25] ), .QN(\mreg/_05074_ ) );
DFF_X1 \mreg/_11684_ ( .CK(clk ), .D(\mreg/_06823_ ), .Q(\mreg/rf[27][26] ), .QN(\mreg/_05073_ ) );
DFF_X1 \mreg/_11685_ ( .CK(clk ), .D(\mreg/_06824_ ), .Q(\mreg/rf[27][27] ), .QN(\mreg/_05072_ ) );
DFF_X1 \mreg/_11686_ ( .CK(clk ), .D(\mreg/_06825_ ), .Q(\mreg/rf[27][28] ), .QN(\mreg/_05071_ ) );
DFF_X1 \mreg/_11687_ ( .CK(clk ), .D(\mreg/_06826_ ), .Q(\mreg/rf[27][29] ), .QN(\mreg/_05070_ ) );
DFF_X1 \mreg/_11688_ ( .CK(clk ), .D(\mreg/_06827_ ), .Q(\mreg/rf[27][30] ), .QN(\mreg/_05069_ ) );
DFF_X1 \mreg/_11689_ ( .CK(clk ), .D(\mreg/_06828_ ), .Q(\mreg/rf[27][31] ), .QN(\mreg/_05068_ ) );
DFF_X1 \mreg/_11690_ ( .CK(clk ), .D(\mreg/_06829_ ), .Q(\mreg/rf[28][0] ), .QN(\mreg/_05067_ ) );
DFF_X1 \mreg/_11691_ ( .CK(clk ), .D(\mreg/_06830_ ), .Q(\mreg/rf[28][1] ), .QN(\mreg/_05066_ ) );
DFF_X1 \mreg/_11692_ ( .CK(clk ), .D(\mreg/_06831_ ), .Q(\mreg/rf[28][2] ), .QN(\mreg/_05065_ ) );
DFF_X1 \mreg/_11693_ ( .CK(clk ), .D(\mreg/_06832_ ), .Q(\mreg/rf[28][3] ), .QN(\mreg/_05064_ ) );
DFF_X1 \mreg/_11694_ ( .CK(clk ), .D(\mreg/_06833_ ), .Q(\mreg/rf[28][4] ), .QN(\mreg/_05063_ ) );
DFF_X1 \mreg/_11695_ ( .CK(clk ), .D(\mreg/_06834_ ), .Q(\mreg/rf[28][5] ), .QN(\mreg/_05062_ ) );
DFF_X1 \mreg/_11696_ ( .CK(clk ), .D(\mreg/_06835_ ), .Q(\mreg/rf[28][6] ), .QN(\mreg/_05061_ ) );
DFF_X1 \mreg/_11697_ ( .CK(clk ), .D(\mreg/_06836_ ), .Q(\mreg/rf[28][7] ), .QN(\mreg/_05060_ ) );
DFF_X1 \mreg/_11698_ ( .CK(clk ), .D(\mreg/_06837_ ), .Q(\mreg/rf[28][8] ), .QN(\mreg/_05059_ ) );
DFF_X1 \mreg/_11699_ ( .CK(clk ), .D(\mreg/_06838_ ), .Q(\mreg/rf[28][9] ), .QN(\mreg/_05058_ ) );
DFF_X1 \mreg/_11700_ ( .CK(clk ), .D(\mreg/_06839_ ), .Q(\mreg/rf[28][10] ), .QN(\mreg/_05057_ ) );
DFF_X1 \mreg/_11701_ ( .CK(clk ), .D(\mreg/_06840_ ), .Q(\mreg/rf[28][11] ), .QN(\mreg/_05056_ ) );
DFF_X1 \mreg/_11702_ ( .CK(clk ), .D(\mreg/_06841_ ), .Q(\mreg/rf[28][12] ), .QN(\mreg/_05055_ ) );
DFF_X1 \mreg/_11703_ ( .CK(clk ), .D(\mreg/_06842_ ), .Q(\mreg/rf[28][13] ), .QN(\mreg/_05054_ ) );
DFF_X1 \mreg/_11704_ ( .CK(clk ), .D(\mreg/_06843_ ), .Q(\mreg/rf[28][14] ), .QN(\mreg/_05053_ ) );
DFF_X1 \mreg/_11705_ ( .CK(clk ), .D(\mreg/_06844_ ), .Q(\mreg/rf[28][15] ), .QN(\mreg/_05052_ ) );
DFF_X1 \mreg/_11706_ ( .CK(clk ), .D(\mreg/_06845_ ), .Q(\mreg/rf[28][16] ), .QN(\mreg/_05051_ ) );
DFF_X1 \mreg/_11707_ ( .CK(clk ), .D(\mreg/_06846_ ), .Q(\mreg/rf[28][17] ), .QN(\mreg/_05050_ ) );
DFF_X1 \mreg/_11708_ ( .CK(clk ), .D(\mreg/_06847_ ), .Q(\mreg/rf[28][18] ), .QN(\mreg/_05049_ ) );
DFF_X1 \mreg/_11709_ ( .CK(clk ), .D(\mreg/_06848_ ), .Q(\mreg/rf[28][19] ), .QN(\mreg/_05048_ ) );
DFF_X1 \mreg/_11710_ ( .CK(clk ), .D(\mreg/_06849_ ), .Q(\mreg/rf[28][20] ), .QN(\mreg/_05047_ ) );
DFF_X1 \mreg/_11711_ ( .CK(clk ), .D(\mreg/_06850_ ), .Q(\mreg/rf[28][21] ), .QN(\mreg/_05046_ ) );
DFF_X1 \mreg/_11712_ ( .CK(clk ), .D(\mreg/_06851_ ), .Q(\mreg/rf[28][22] ), .QN(\mreg/_05045_ ) );
DFF_X1 \mreg/_11713_ ( .CK(clk ), .D(\mreg/_06852_ ), .Q(\mreg/rf[28][23] ), .QN(\mreg/_05044_ ) );
DFF_X1 \mreg/_11714_ ( .CK(clk ), .D(\mreg/_06853_ ), .Q(\mreg/rf[28][24] ), .QN(\mreg/_05043_ ) );
DFF_X1 \mreg/_11715_ ( .CK(clk ), .D(\mreg/_06854_ ), .Q(\mreg/rf[28][25] ), .QN(\mreg/_05042_ ) );
DFF_X1 \mreg/_11716_ ( .CK(clk ), .D(\mreg/_06855_ ), .Q(\mreg/rf[28][26] ), .QN(\mreg/_05041_ ) );
DFF_X1 \mreg/_11717_ ( .CK(clk ), .D(\mreg/_06856_ ), .Q(\mreg/rf[28][27] ), .QN(\mreg/_05040_ ) );
DFF_X1 \mreg/_11718_ ( .CK(clk ), .D(\mreg/_06857_ ), .Q(\mreg/rf[28][28] ), .QN(\mreg/_05039_ ) );
DFF_X1 \mreg/_11719_ ( .CK(clk ), .D(\mreg/_06858_ ), .Q(\mreg/rf[28][29] ), .QN(\mreg/_05038_ ) );
DFF_X1 \mreg/_11720_ ( .CK(clk ), .D(\mreg/_06859_ ), .Q(\mreg/rf[28][30] ), .QN(\mreg/_05037_ ) );
DFF_X1 \mreg/_11721_ ( .CK(clk ), .D(\mreg/_06860_ ), .Q(\mreg/rf[28][31] ), .QN(\mreg/_05036_ ) );
DFF_X1 \mreg/_11722_ ( .CK(clk ), .D(\mreg/_06861_ ), .Q(\mreg/rf[29][0] ), .QN(\mreg/_05035_ ) );
DFF_X1 \mreg/_11723_ ( .CK(clk ), .D(\mreg/_06862_ ), .Q(\mreg/rf[29][1] ), .QN(\mreg/_05034_ ) );
DFF_X1 \mreg/_11724_ ( .CK(clk ), .D(\mreg/_06863_ ), .Q(\mreg/rf[29][2] ), .QN(\mreg/_05033_ ) );
DFF_X1 \mreg/_11725_ ( .CK(clk ), .D(\mreg/_06864_ ), .Q(\mreg/rf[29][3] ), .QN(\mreg/_05032_ ) );
DFF_X1 \mreg/_11726_ ( .CK(clk ), .D(\mreg/_06865_ ), .Q(\mreg/rf[29][4] ), .QN(\mreg/_05031_ ) );
DFF_X1 \mreg/_11727_ ( .CK(clk ), .D(\mreg/_06866_ ), .Q(\mreg/rf[29][5] ), .QN(\mreg/_05030_ ) );
DFF_X1 \mreg/_11728_ ( .CK(clk ), .D(\mreg/_06867_ ), .Q(\mreg/rf[29][6] ), .QN(\mreg/_05029_ ) );
DFF_X1 \mreg/_11729_ ( .CK(clk ), .D(\mreg/_06868_ ), .Q(\mreg/rf[29][7] ), .QN(\mreg/_05028_ ) );
DFF_X1 \mreg/_11730_ ( .CK(clk ), .D(\mreg/_06869_ ), .Q(\mreg/rf[29][8] ), .QN(\mreg/_05027_ ) );
DFF_X1 \mreg/_11731_ ( .CK(clk ), .D(\mreg/_06870_ ), .Q(\mreg/rf[29][9] ), .QN(\mreg/_05026_ ) );
DFF_X1 \mreg/_11732_ ( .CK(clk ), .D(\mreg/_06871_ ), .Q(\mreg/rf[29][10] ), .QN(\mreg/_05025_ ) );
DFF_X1 \mreg/_11733_ ( .CK(clk ), .D(\mreg/_06872_ ), .Q(\mreg/rf[29][11] ), .QN(\mreg/_05024_ ) );
DFF_X1 \mreg/_11734_ ( .CK(clk ), .D(\mreg/_06873_ ), .Q(\mreg/rf[29][12] ), .QN(\mreg/_05023_ ) );
DFF_X1 \mreg/_11735_ ( .CK(clk ), .D(\mreg/_06874_ ), .Q(\mreg/rf[29][13] ), .QN(\mreg/_05022_ ) );
DFF_X1 \mreg/_11736_ ( .CK(clk ), .D(\mreg/_06875_ ), .Q(\mreg/rf[29][14] ), .QN(\mreg/_05021_ ) );
DFF_X1 \mreg/_11737_ ( .CK(clk ), .D(\mreg/_06876_ ), .Q(\mreg/rf[29][15] ), .QN(\mreg/_05020_ ) );
DFF_X1 \mreg/_11738_ ( .CK(clk ), .D(\mreg/_06877_ ), .Q(\mreg/rf[29][16] ), .QN(\mreg/_05019_ ) );
DFF_X1 \mreg/_11739_ ( .CK(clk ), .D(\mreg/_06878_ ), .Q(\mreg/rf[29][17] ), .QN(\mreg/_05018_ ) );
DFF_X1 \mreg/_11740_ ( .CK(clk ), .D(\mreg/_06879_ ), .Q(\mreg/rf[29][18] ), .QN(\mreg/_05017_ ) );
DFF_X1 \mreg/_11741_ ( .CK(clk ), .D(\mreg/_06880_ ), .Q(\mreg/rf[29][19] ), .QN(\mreg/_05016_ ) );
DFF_X1 \mreg/_11742_ ( .CK(clk ), .D(\mreg/_06881_ ), .Q(\mreg/rf[29][20] ), .QN(\mreg/_05015_ ) );
DFF_X1 \mreg/_11743_ ( .CK(clk ), .D(\mreg/_06882_ ), .Q(\mreg/rf[29][21] ), .QN(\mreg/_05014_ ) );
DFF_X1 \mreg/_11744_ ( .CK(clk ), .D(\mreg/_06883_ ), .Q(\mreg/rf[29][22] ), .QN(\mreg/_05013_ ) );
DFF_X1 \mreg/_11745_ ( .CK(clk ), .D(\mreg/_06884_ ), .Q(\mreg/rf[29][23] ), .QN(\mreg/_05012_ ) );
DFF_X1 \mreg/_11746_ ( .CK(clk ), .D(\mreg/_06885_ ), .Q(\mreg/rf[29][24] ), .QN(\mreg/_05011_ ) );
DFF_X1 \mreg/_11747_ ( .CK(clk ), .D(\mreg/_06886_ ), .Q(\mreg/rf[29][25] ), .QN(\mreg/_05010_ ) );
DFF_X1 \mreg/_11748_ ( .CK(clk ), .D(\mreg/_06887_ ), .Q(\mreg/rf[29][26] ), .QN(\mreg/_05009_ ) );
DFF_X1 \mreg/_11749_ ( .CK(clk ), .D(\mreg/_06888_ ), .Q(\mreg/rf[29][27] ), .QN(\mreg/_05008_ ) );
DFF_X1 \mreg/_11750_ ( .CK(clk ), .D(\mreg/_06889_ ), .Q(\mreg/rf[29][28] ), .QN(\mreg/_05007_ ) );
DFF_X1 \mreg/_11751_ ( .CK(clk ), .D(\mreg/_06890_ ), .Q(\mreg/rf[29][29] ), .QN(\mreg/_05006_ ) );
DFF_X1 \mreg/_11752_ ( .CK(clk ), .D(\mreg/_06891_ ), .Q(\mreg/rf[29][30] ), .QN(\mreg/_05005_ ) );
DFF_X1 \mreg/_11753_ ( .CK(clk ), .D(\mreg/_06892_ ), .Q(\mreg/rf[29][31] ), .QN(\mreg/_05004_ ) );
DFF_X1 \mreg/_11754_ ( .CK(clk ), .D(\mreg/_06893_ ), .Q(\mreg/rf[30][0] ), .QN(\mreg/_05003_ ) );
DFF_X1 \mreg/_11755_ ( .CK(clk ), .D(\mreg/_06894_ ), .Q(\mreg/rf[30][1] ), .QN(\mreg/_05002_ ) );
DFF_X1 \mreg/_11756_ ( .CK(clk ), .D(\mreg/_06895_ ), .Q(\mreg/rf[30][2] ), .QN(\mreg/_05001_ ) );
DFF_X1 \mreg/_11757_ ( .CK(clk ), .D(\mreg/_06896_ ), .Q(\mreg/rf[30][3] ), .QN(\mreg/_05000_ ) );
DFF_X1 \mreg/_11758_ ( .CK(clk ), .D(\mreg/_06897_ ), .Q(\mreg/rf[30][4] ), .QN(\mreg/_04999_ ) );
DFF_X1 \mreg/_11759_ ( .CK(clk ), .D(\mreg/_06898_ ), .Q(\mreg/rf[30][5] ), .QN(\mreg/_04998_ ) );
DFF_X1 \mreg/_11760_ ( .CK(clk ), .D(\mreg/_06899_ ), .Q(\mreg/rf[30][6] ), .QN(\mreg/_04997_ ) );
DFF_X1 \mreg/_11761_ ( .CK(clk ), .D(\mreg/_06900_ ), .Q(\mreg/rf[30][7] ), .QN(\mreg/_04996_ ) );
DFF_X1 \mreg/_11762_ ( .CK(clk ), .D(\mreg/_06901_ ), .Q(\mreg/rf[30][8] ), .QN(\mreg/_04995_ ) );
DFF_X1 \mreg/_11763_ ( .CK(clk ), .D(\mreg/_06902_ ), .Q(\mreg/rf[30][9] ), .QN(\mreg/_04994_ ) );
DFF_X1 \mreg/_11764_ ( .CK(clk ), .D(\mreg/_06903_ ), .Q(\mreg/rf[30][10] ), .QN(\mreg/_04993_ ) );
DFF_X1 \mreg/_11765_ ( .CK(clk ), .D(\mreg/_06904_ ), .Q(\mreg/rf[30][11] ), .QN(\mreg/_04992_ ) );
DFF_X1 \mreg/_11766_ ( .CK(clk ), .D(\mreg/_06905_ ), .Q(\mreg/rf[30][12] ), .QN(\mreg/_04991_ ) );
DFF_X1 \mreg/_11767_ ( .CK(clk ), .D(\mreg/_06906_ ), .Q(\mreg/rf[30][13] ), .QN(\mreg/_04990_ ) );
DFF_X1 \mreg/_11768_ ( .CK(clk ), .D(\mreg/_06907_ ), .Q(\mreg/rf[30][14] ), .QN(\mreg/_04989_ ) );
DFF_X1 \mreg/_11769_ ( .CK(clk ), .D(\mreg/_06908_ ), .Q(\mreg/rf[30][15] ), .QN(\mreg/_04988_ ) );
DFF_X1 \mreg/_11770_ ( .CK(clk ), .D(\mreg/_06909_ ), .Q(\mreg/rf[30][16] ), .QN(\mreg/_04987_ ) );
DFF_X1 \mreg/_11771_ ( .CK(clk ), .D(\mreg/_06910_ ), .Q(\mreg/rf[30][17] ), .QN(\mreg/_04986_ ) );
DFF_X1 \mreg/_11772_ ( .CK(clk ), .D(\mreg/_06911_ ), .Q(\mreg/rf[30][18] ), .QN(\mreg/_04985_ ) );
DFF_X1 \mreg/_11773_ ( .CK(clk ), .D(\mreg/_06912_ ), .Q(\mreg/rf[30][19] ), .QN(\mreg/_04984_ ) );
DFF_X1 \mreg/_11774_ ( .CK(clk ), .D(\mreg/_06913_ ), .Q(\mreg/rf[30][20] ), .QN(\mreg/_04983_ ) );
DFF_X1 \mreg/_11775_ ( .CK(clk ), .D(\mreg/_06914_ ), .Q(\mreg/rf[30][21] ), .QN(\mreg/_04982_ ) );
DFF_X1 \mreg/_11776_ ( .CK(clk ), .D(\mreg/_06915_ ), .Q(\mreg/rf[30][22] ), .QN(\mreg/_04981_ ) );
DFF_X1 \mreg/_11777_ ( .CK(clk ), .D(\mreg/_06916_ ), .Q(\mreg/rf[30][23] ), .QN(\mreg/_04980_ ) );
DFF_X1 \mreg/_11778_ ( .CK(clk ), .D(\mreg/_06917_ ), .Q(\mreg/rf[30][24] ), .QN(\mreg/_04979_ ) );
DFF_X1 \mreg/_11779_ ( .CK(clk ), .D(\mreg/_06918_ ), .Q(\mreg/rf[30][25] ), .QN(\mreg/_04978_ ) );
DFF_X1 \mreg/_11780_ ( .CK(clk ), .D(\mreg/_06919_ ), .Q(\mreg/rf[30][26] ), .QN(\mreg/_04977_ ) );
DFF_X1 \mreg/_11781_ ( .CK(clk ), .D(\mreg/_06920_ ), .Q(\mreg/rf[30][27] ), .QN(\mreg/_04976_ ) );
DFF_X1 \mreg/_11782_ ( .CK(clk ), .D(\mreg/_06921_ ), .Q(\mreg/rf[30][28] ), .QN(\mreg/_04975_ ) );
DFF_X1 \mreg/_11783_ ( .CK(clk ), .D(\mreg/_06922_ ), .Q(\mreg/rf[30][29] ), .QN(\mreg/_04974_ ) );
DFF_X1 \mreg/_11784_ ( .CK(clk ), .D(\mreg/_06923_ ), .Q(\mreg/rf[30][30] ), .QN(\mreg/_04973_ ) );
DFF_X1 \mreg/_11785_ ( .CK(clk ), .D(\mreg/_06924_ ), .Q(\mreg/rf[30][31] ), .QN(\mreg/_04972_ ) );
BUF_X1 \mreg/_11786_ ( .A(reg_wen ), .Z(\mreg/_04971_ ) );
BUF_X1 \mreg/_11787_ ( .A(lsu_finish ), .Z(\mreg/_01054_ ) );
BUF_X1 \mreg/_11788_ ( .A(\rd[4] ), .Z(\mreg/_04938_ ) );
BUF_X1 \mreg/_11789_ ( .A(\rd[0] ), .Z(\mreg/_04934_ ) );
BUF_X1 \mreg/_11790_ ( .A(\rd[1] ), .Z(\mreg/_04935_ ) );
BUF_X1 \mreg/_11791_ ( .A(\rd[2] ), .Z(\mreg/_04936_ ) );
BUF_X1 \mreg/_11792_ ( .A(\rd[3] ), .Z(\mreg/_04937_ ) );
BUF_X1 \mreg/_11793_ ( .A(\rs2[4] ), .Z(\mreg/_03877_ ) );
BUF_X1 \mreg/_11794_ ( .A(\rs2[1] ), .Z(\mreg/_03874_ ) );
BUF_X1 \mreg/_11795_ ( .A(\rs2[0] ), .Z(\mreg/_03873_ ) );
BUF_X1 \mreg/_11796_ ( .A(\rs2[3] ), .Z(\mreg/_03876_ ) );
BUF_X1 \mreg/_11797_ ( .A(\rs2[2] ), .Z(\mreg/_03875_ ) );
BUF_X1 \mreg/_11798_ ( .A(\mreg/rf[31][0] ), .Z(\mreg/_04678_ ) );
BUF_X1 \mreg/_11799_ ( .A(\mreg/rf[30][0] ), .Z(\mreg/_04646_ ) );
BUF_X1 \mreg/_11800_ ( .A(\mreg/rf[29][0] ), .Z(\mreg/_04582_ ) );
BUF_X1 \mreg/_11801_ ( .A(\mreg/rf[28][0] ), .Z(\mreg/_04550_ ) );
BUF_X1 \mreg/_11802_ ( .A(\mreg/rf[27][0] ), .Z(\mreg/_04518_ ) );
BUF_X1 \mreg/_11803_ ( .A(\mreg/rf[26][0] ), .Z(\mreg/_04486_ ) );
BUF_X1 \mreg/_11804_ ( .A(\mreg/rf[25][0] ), .Z(\mreg/_04454_ ) );
BUF_X1 \mreg/_11805_ ( .A(\mreg/rf[24][0] ), .Z(\mreg/_04422_ ) );
BUF_X1 \mreg/_11806_ ( .A(\mreg/rf[23][0] ), .Z(\mreg/_04390_ ) );
BUF_X1 \mreg/_11807_ ( .A(\mreg/rf[22][0] ), .Z(\mreg/_04358_ ) );
BUF_X1 \mreg/_11808_ ( .A(\mreg/rf[21][0] ), .Z(\mreg/_04326_ ) );
BUF_X1 \mreg/_11809_ ( .A(\mreg/rf[20][0] ), .Z(\mreg/_04294_ ) );
BUF_X1 \mreg/_11810_ ( .A(\mreg/rf[19][0] ), .Z(\mreg/_04230_ ) );
BUF_X1 \mreg/_11811_ ( .A(\mreg/rf[18][0] ), .Z(\mreg/_04198_ ) );
BUF_X1 \mreg/_11812_ ( .A(\mreg/rf[17][0] ), .Z(\mreg/_04166_ ) );
BUF_X1 \mreg/_11813_ ( .A(\mreg/rf[16][0] ), .Z(\mreg/_04134_ ) );
BUF_X1 \mreg/_11814_ ( .A(\mreg/rf[15][0] ), .Z(\mreg/_04102_ ) );
BUF_X1 \mreg/_11815_ ( .A(\mreg/rf[14][0] ), .Z(\mreg/_04070_ ) );
BUF_X1 \mreg/_11816_ ( .A(\mreg/rf[13][0] ), .Z(\mreg/_04038_ ) );
BUF_X1 \mreg/_11817_ ( .A(\mreg/rf[12][0] ), .Z(\mreg/_04006_ ) );
BUF_X1 \mreg/_11818_ ( .A(\mreg/rf[11][0] ), .Z(\mreg/_03974_ ) );
BUF_X1 \mreg/_11819_ ( .A(\mreg/rf[10][0] ), .Z(\mreg/_03942_ ) );
BUF_X1 \mreg/_11820_ ( .A(\mreg/rf[9][0] ), .Z(\mreg/_04902_ ) );
BUF_X1 \mreg/_11821_ ( .A(\mreg/rf[8][0] ), .Z(\mreg/_04870_ ) );
BUF_X1 \mreg/_11822_ ( .A(\mreg/rf[7][0] ), .Z(\mreg/_04838_ ) );
BUF_X1 \mreg/_11823_ ( .A(\mreg/rf[6][0] ), .Z(\mreg/_04806_ ) );
BUF_X1 \mreg/_11824_ ( .A(\mreg/rf[5][0] ), .Z(\mreg/_04774_ ) );
BUF_X1 \mreg/_11825_ ( .A(\mreg/rf[4][0] ), .Z(\mreg/_04742_ ) );
BUF_X1 \mreg/_11826_ ( .A(\mreg/rf[3][0] ), .Z(\mreg/_04710_ ) );
BUF_X1 \mreg/_11827_ ( .A(\mreg/rf[2][0] ), .Z(\mreg/_04614_ ) );
BUF_X1 \mreg/_11828_ ( .A(\mreg/rf[1][0] ), .Z(\mreg/_04262_ ) );
BUF_X1 \mreg/_11829_ ( .A(\mreg/_03910_ ), .Z(\mem_wdata[0] ) );
BUF_X1 \mreg/_11830_ ( .A(\mreg/_00000_ ), .Z(\mreg/_00031_ ) );
BUF_X1 \mreg/_11831_ ( .A(\mreg/rf[30][1] ), .Z(\mreg/_04657_ ) );
BUF_X1 \mreg/_11832_ ( .A(\mreg/rf[29][1] ), .Z(\mreg/_04593_ ) );
BUF_X1 \mreg/_11833_ ( .A(\mreg/rf[28][1] ), .Z(\mreg/_04561_ ) );
BUF_X1 \mreg/_11834_ ( .A(\mreg/rf[27][1] ), .Z(\mreg/_04529_ ) );
BUF_X1 \mreg/_11835_ ( .A(\mreg/rf[26][1] ), .Z(\mreg/_04497_ ) );
BUF_X1 \mreg/_11836_ ( .A(\mreg/rf[25][1] ), .Z(\mreg/_04465_ ) );
BUF_X1 \mreg/_11837_ ( .A(\mreg/rf[24][1] ), .Z(\mreg/_04433_ ) );
BUF_X1 \mreg/_11838_ ( .A(\mreg/rf[23][1] ), .Z(\mreg/_04401_ ) );
BUF_X1 \mreg/_11839_ ( .A(\mreg/rf[22][1] ), .Z(\mreg/_04369_ ) );
BUF_X1 \mreg/_11840_ ( .A(\mreg/rf[21][1] ), .Z(\mreg/_04337_ ) );
BUF_X1 \mreg/_11841_ ( .A(\mreg/rf[20][1] ), .Z(\mreg/_04305_ ) );
BUF_X1 \mreg/_11842_ ( .A(\mreg/rf[19][1] ), .Z(\mreg/_04241_ ) );
BUF_X1 \mreg/_11843_ ( .A(\mreg/rf[18][1] ), .Z(\mreg/_04209_ ) );
BUF_X1 \mreg/_11844_ ( .A(\mreg/rf[17][1] ), .Z(\mreg/_04177_ ) );
BUF_X1 \mreg/_11845_ ( .A(\mreg/rf[16][1] ), .Z(\mreg/_04145_ ) );
BUF_X1 \mreg/_11846_ ( .A(\mreg/rf[15][1] ), .Z(\mreg/_04113_ ) );
BUF_X1 \mreg/_11847_ ( .A(\mreg/rf[14][1] ), .Z(\mreg/_04081_ ) );
BUF_X1 \mreg/_11848_ ( .A(\mreg/rf[13][1] ), .Z(\mreg/_04049_ ) );
BUF_X1 \mreg/_11849_ ( .A(\mreg/rf[12][1] ), .Z(\mreg/_04017_ ) );
BUF_X1 \mreg/_11850_ ( .A(\mreg/rf[11][1] ), .Z(\mreg/_03985_ ) );
BUF_X1 \mreg/_11851_ ( .A(\mreg/rf[10][1] ), .Z(\mreg/_03953_ ) );
BUF_X1 \mreg/_11852_ ( .A(\mreg/rf[9][1] ), .Z(\mreg/_04913_ ) );
BUF_X1 \mreg/_11853_ ( .A(\mreg/rf[8][1] ), .Z(\mreg/_04881_ ) );
BUF_X1 \mreg/_11854_ ( .A(\mreg/rf[7][1] ), .Z(\mreg/_04849_ ) );
BUF_X1 \mreg/_11855_ ( .A(\mreg/rf[6][1] ), .Z(\mreg/_04817_ ) );
BUF_X1 \mreg/_11856_ ( .A(\mreg/rf[5][1] ), .Z(\mreg/_04785_ ) );
BUF_X1 \mreg/_11857_ ( .A(\mreg/rf[4][1] ), .Z(\mreg/_04753_ ) );
BUF_X1 \mreg/_11858_ ( .A(\mreg/rf[3][1] ), .Z(\mreg/_04721_ ) );
BUF_X1 \mreg/_11859_ ( .A(\mreg/rf[2][1] ), .Z(\mreg/_04625_ ) );
BUF_X1 \mreg/_11860_ ( .A(\mreg/rf[1][1] ), .Z(\mreg/_04273_ ) );
BUF_X1 \mreg/_11861_ ( .A(\mreg/_03921_ ), .Z(\mem_wdata[1] ) );
BUF_X1 \mreg/_11862_ ( .A(\mreg/_00001_ ), .Z(\mreg/_00032_ ) );
BUF_X1 \mreg/_11863_ ( .A(\mreg/rf[30][2] ), .Z(\mreg/_04668_ ) );
BUF_X1 \mreg/_11864_ ( .A(\mreg/rf[29][2] ), .Z(\mreg/_04604_ ) );
BUF_X1 \mreg/_11865_ ( .A(\mreg/rf[28][2] ), .Z(\mreg/_04572_ ) );
BUF_X1 \mreg/_11866_ ( .A(\mreg/rf[27][2] ), .Z(\mreg/_04540_ ) );
BUF_X1 \mreg/_11867_ ( .A(\mreg/rf[26][2] ), .Z(\mreg/_04508_ ) );
BUF_X1 \mreg/_11868_ ( .A(\mreg/rf[25][2] ), .Z(\mreg/_04476_ ) );
BUF_X1 \mreg/_11869_ ( .A(\mreg/rf[24][2] ), .Z(\mreg/_04444_ ) );
BUF_X1 \mreg/_11870_ ( .A(\mreg/rf[23][2] ), .Z(\mreg/_04412_ ) );
BUF_X1 \mreg/_11871_ ( .A(\mreg/rf[22][2] ), .Z(\mreg/_04380_ ) );
BUF_X1 \mreg/_11872_ ( .A(\mreg/rf[21][2] ), .Z(\mreg/_04348_ ) );
BUF_X1 \mreg/_11873_ ( .A(\mreg/rf[20][2] ), .Z(\mreg/_04316_ ) );
BUF_X1 \mreg/_11874_ ( .A(\mreg/rf[19][2] ), .Z(\mreg/_04252_ ) );
BUF_X1 \mreg/_11875_ ( .A(\mreg/rf[18][2] ), .Z(\mreg/_04220_ ) );
BUF_X1 \mreg/_11876_ ( .A(\mreg/rf[17][2] ), .Z(\mreg/_04188_ ) );
BUF_X1 \mreg/_11877_ ( .A(\mreg/rf[16][2] ), .Z(\mreg/_04156_ ) );
BUF_X1 \mreg/_11878_ ( .A(\mreg/rf[15][2] ), .Z(\mreg/_04124_ ) );
BUF_X1 \mreg/_11879_ ( .A(\mreg/rf[14][2] ), .Z(\mreg/_04092_ ) );
BUF_X1 \mreg/_11880_ ( .A(\mreg/rf[13][2] ), .Z(\mreg/_04060_ ) );
BUF_X1 \mreg/_11881_ ( .A(\mreg/rf[12][2] ), .Z(\mreg/_04028_ ) );
BUF_X1 \mreg/_11882_ ( .A(\mreg/rf[11][2] ), .Z(\mreg/_03996_ ) );
BUF_X1 \mreg/_11883_ ( .A(\mreg/rf[10][2] ), .Z(\mreg/_03964_ ) );
BUF_X1 \mreg/_11884_ ( .A(\mreg/rf[9][2] ), .Z(\mreg/_04924_ ) );
BUF_X1 \mreg/_11885_ ( .A(\mreg/rf[8][2] ), .Z(\mreg/_04892_ ) );
BUF_X1 \mreg/_11886_ ( .A(\mreg/rf[7][2] ), .Z(\mreg/_04860_ ) );
BUF_X1 \mreg/_11887_ ( .A(\mreg/rf[6][2] ), .Z(\mreg/_04828_ ) );
BUF_X1 \mreg/_11888_ ( .A(\mreg/rf[5][2] ), .Z(\mreg/_04796_ ) );
BUF_X1 \mreg/_11889_ ( .A(\mreg/rf[4][2] ), .Z(\mreg/_04764_ ) );
BUF_X1 \mreg/_11890_ ( .A(\mreg/rf[3][2] ), .Z(\mreg/_04732_ ) );
BUF_X1 \mreg/_11891_ ( .A(\mreg/rf[2][2] ), .Z(\mreg/_04636_ ) );
BUF_X1 \mreg/_11892_ ( .A(\mreg/rf[1][2] ), .Z(\mreg/_04284_ ) );
BUF_X1 \mreg/_11893_ ( .A(\mreg/_03932_ ), .Z(\mem_wdata[2] ) );
BUF_X1 \mreg/_11894_ ( .A(\mreg/_00002_ ), .Z(\mreg/_00033_ ) );
BUF_X1 \mreg/_11895_ ( .A(\mreg/rf[30][3] ), .Z(\mreg/_04671_ ) );
BUF_X1 \mreg/_11896_ ( .A(\mreg/rf[29][3] ), .Z(\mreg/_04607_ ) );
BUF_X1 \mreg/_11897_ ( .A(\mreg/rf[28][3] ), .Z(\mreg/_04575_ ) );
BUF_X1 \mreg/_11898_ ( .A(\mreg/rf[27][3] ), .Z(\mreg/_04543_ ) );
BUF_X1 \mreg/_11899_ ( .A(\mreg/rf[26][3] ), .Z(\mreg/_04511_ ) );
BUF_X1 \mreg/_11900_ ( .A(\mreg/rf[25][3] ), .Z(\mreg/_04479_ ) );
BUF_X1 \mreg/_11901_ ( .A(\mreg/rf[24][3] ), .Z(\mreg/_04447_ ) );
BUF_X1 \mreg/_11902_ ( .A(\mreg/rf[23][3] ), .Z(\mreg/_04415_ ) );
BUF_X1 \mreg/_11903_ ( .A(\mreg/rf[22][3] ), .Z(\mreg/_04383_ ) );
BUF_X1 \mreg/_11904_ ( .A(\mreg/rf[21][3] ), .Z(\mreg/_04351_ ) );
BUF_X1 \mreg/_11905_ ( .A(\mreg/rf[20][3] ), .Z(\mreg/_04319_ ) );
BUF_X1 \mreg/_11906_ ( .A(\mreg/rf[19][3] ), .Z(\mreg/_04255_ ) );
BUF_X1 \mreg/_11907_ ( .A(\mreg/rf[18][3] ), .Z(\mreg/_04223_ ) );
BUF_X1 \mreg/_11908_ ( .A(\mreg/rf[17][3] ), .Z(\mreg/_04191_ ) );
BUF_X1 \mreg/_11909_ ( .A(\mreg/rf[16][3] ), .Z(\mreg/_04159_ ) );
BUF_X1 \mreg/_11910_ ( .A(\mreg/rf[15][3] ), .Z(\mreg/_04127_ ) );
BUF_X1 \mreg/_11911_ ( .A(\mreg/rf[14][3] ), .Z(\mreg/_04095_ ) );
BUF_X1 \mreg/_11912_ ( .A(\mreg/rf[13][3] ), .Z(\mreg/_04063_ ) );
BUF_X1 \mreg/_11913_ ( .A(\mreg/rf[12][3] ), .Z(\mreg/_04031_ ) );
BUF_X1 \mreg/_11914_ ( .A(\mreg/rf[11][3] ), .Z(\mreg/_03999_ ) );
BUF_X1 \mreg/_11915_ ( .A(\mreg/rf[10][3] ), .Z(\mreg/_03967_ ) );
BUF_X1 \mreg/_11916_ ( .A(\mreg/rf[9][3] ), .Z(\mreg/_04927_ ) );
BUF_X1 \mreg/_11917_ ( .A(\mreg/rf[8][3] ), .Z(\mreg/_04895_ ) );
BUF_X1 \mreg/_11918_ ( .A(\mreg/rf[7][3] ), .Z(\mreg/_04863_ ) );
BUF_X1 \mreg/_11919_ ( .A(\mreg/rf[6][3] ), .Z(\mreg/_04831_ ) );
BUF_X1 \mreg/_11920_ ( .A(\mreg/rf[5][3] ), .Z(\mreg/_04799_ ) );
BUF_X1 \mreg/_11921_ ( .A(\mreg/rf[4][3] ), .Z(\mreg/_04767_ ) );
BUF_X1 \mreg/_11922_ ( .A(\mreg/rf[3][3] ), .Z(\mreg/_04735_ ) );
BUF_X1 \mreg/_11923_ ( .A(\mreg/rf[2][3] ), .Z(\mreg/_04639_ ) );
BUF_X1 \mreg/_11924_ ( .A(\mreg/rf[1][3] ), .Z(\mreg/_04287_ ) );
BUF_X1 \mreg/_11925_ ( .A(\mreg/_03935_ ), .Z(\mem_wdata[3] ) );
BUF_X1 \mreg/_11926_ ( .A(\mreg/_00003_ ), .Z(\mreg/_00034_ ) );
BUF_X1 \mreg/_11927_ ( .A(\mreg/rf[30][4] ), .Z(\mreg/_04672_ ) );
BUF_X1 \mreg/_11928_ ( .A(\mreg/rf[29][4] ), .Z(\mreg/_04608_ ) );
BUF_X1 \mreg/_11929_ ( .A(\mreg/rf[28][4] ), .Z(\mreg/_04576_ ) );
BUF_X1 \mreg/_11930_ ( .A(\mreg/rf[27][4] ), .Z(\mreg/_04544_ ) );
BUF_X1 \mreg/_11931_ ( .A(\mreg/rf[26][4] ), .Z(\mreg/_04512_ ) );
BUF_X1 \mreg/_11932_ ( .A(\mreg/rf[25][4] ), .Z(\mreg/_04480_ ) );
BUF_X1 \mreg/_11933_ ( .A(\mreg/rf[24][4] ), .Z(\mreg/_04448_ ) );
BUF_X1 \mreg/_11934_ ( .A(\mreg/rf[23][4] ), .Z(\mreg/_04416_ ) );
BUF_X1 \mreg/_11935_ ( .A(\mreg/rf[22][4] ), .Z(\mreg/_04384_ ) );
BUF_X1 \mreg/_11936_ ( .A(\mreg/rf[21][4] ), .Z(\mreg/_04352_ ) );
BUF_X1 \mreg/_11937_ ( .A(\mreg/rf[20][4] ), .Z(\mreg/_04320_ ) );
BUF_X1 \mreg/_11938_ ( .A(\mreg/rf[19][4] ), .Z(\mreg/_04256_ ) );
BUF_X1 \mreg/_11939_ ( .A(\mreg/rf[18][4] ), .Z(\mreg/_04224_ ) );
BUF_X1 \mreg/_11940_ ( .A(\mreg/rf[17][4] ), .Z(\mreg/_04192_ ) );
BUF_X1 \mreg/_11941_ ( .A(\mreg/rf[16][4] ), .Z(\mreg/_04160_ ) );
BUF_X1 \mreg/_11942_ ( .A(\mreg/rf[15][4] ), .Z(\mreg/_04128_ ) );
BUF_X1 \mreg/_11943_ ( .A(\mreg/rf[14][4] ), .Z(\mreg/_04096_ ) );
BUF_X1 \mreg/_11944_ ( .A(\mreg/rf[13][4] ), .Z(\mreg/_04064_ ) );
BUF_X1 \mreg/_11945_ ( .A(\mreg/rf[12][4] ), .Z(\mreg/_04032_ ) );
BUF_X1 \mreg/_11946_ ( .A(\mreg/rf[11][4] ), .Z(\mreg/_04000_ ) );
BUF_X1 \mreg/_11947_ ( .A(\mreg/rf[10][4] ), .Z(\mreg/_03968_ ) );
BUF_X1 \mreg/_11948_ ( .A(\mreg/rf[9][4] ), .Z(\mreg/_04928_ ) );
BUF_X1 \mreg/_11949_ ( .A(\mreg/rf[8][4] ), .Z(\mreg/_04896_ ) );
BUF_X1 \mreg/_11950_ ( .A(\mreg/rf[7][4] ), .Z(\mreg/_04864_ ) );
BUF_X1 \mreg/_11951_ ( .A(\mreg/rf[6][4] ), .Z(\mreg/_04832_ ) );
BUF_X1 \mreg/_11952_ ( .A(\mreg/rf[5][4] ), .Z(\mreg/_04800_ ) );
BUF_X1 \mreg/_11953_ ( .A(\mreg/rf[4][4] ), .Z(\mreg/_04768_ ) );
BUF_X1 \mreg/_11954_ ( .A(\mreg/rf[3][4] ), .Z(\mreg/_04736_ ) );
BUF_X1 \mreg/_11955_ ( .A(\mreg/rf[2][4] ), .Z(\mreg/_04640_ ) );
BUF_X1 \mreg/_11956_ ( .A(\mreg/rf[1][4] ), .Z(\mreg/_04288_ ) );
BUF_X1 \mreg/_11957_ ( .A(\mreg/_03936_ ), .Z(\mem_wdata[4] ) );
BUF_X1 \mreg/_11958_ ( .A(\mreg/_00004_ ), .Z(\mreg/_00035_ ) );
BUF_X1 \mreg/_11959_ ( .A(\mreg/rf[30][5] ), .Z(\mreg/_04673_ ) );
BUF_X1 \mreg/_11960_ ( .A(\mreg/rf[29][5] ), .Z(\mreg/_04609_ ) );
BUF_X1 \mreg/_11961_ ( .A(\mreg/rf[28][5] ), .Z(\mreg/_04577_ ) );
BUF_X1 \mreg/_11962_ ( .A(\mreg/rf[27][5] ), .Z(\mreg/_04545_ ) );
BUF_X1 \mreg/_11963_ ( .A(\mreg/rf[26][5] ), .Z(\mreg/_04513_ ) );
BUF_X1 \mreg/_11964_ ( .A(\mreg/rf[25][5] ), .Z(\mreg/_04481_ ) );
BUF_X1 \mreg/_11965_ ( .A(\mreg/rf[24][5] ), .Z(\mreg/_04449_ ) );
BUF_X1 \mreg/_11966_ ( .A(\mreg/rf[23][5] ), .Z(\mreg/_04417_ ) );
BUF_X1 \mreg/_11967_ ( .A(\mreg/rf[22][5] ), .Z(\mreg/_04385_ ) );
BUF_X1 \mreg/_11968_ ( .A(\mreg/rf[21][5] ), .Z(\mreg/_04353_ ) );
BUF_X1 \mreg/_11969_ ( .A(\mreg/rf[20][5] ), .Z(\mreg/_04321_ ) );
BUF_X1 \mreg/_11970_ ( .A(\mreg/rf[19][5] ), .Z(\mreg/_04257_ ) );
BUF_X1 \mreg/_11971_ ( .A(\mreg/rf[18][5] ), .Z(\mreg/_04225_ ) );
BUF_X1 \mreg/_11972_ ( .A(\mreg/rf[17][5] ), .Z(\mreg/_04193_ ) );
BUF_X1 \mreg/_11973_ ( .A(\mreg/rf[16][5] ), .Z(\mreg/_04161_ ) );
BUF_X1 \mreg/_11974_ ( .A(\mreg/rf[15][5] ), .Z(\mreg/_04129_ ) );
BUF_X1 \mreg/_11975_ ( .A(\mreg/rf[14][5] ), .Z(\mreg/_04097_ ) );
BUF_X1 \mreg/_11976_ ( .A(\mreg/rf[13][5] ), .Z(\mreg/_04065_ ) );
BUF_X1 \mreg/_11977_ ( .A(\mreg/rf[12][5] ), .Z(\mreg/_04033_ ) );
BUF_X1 \mreg/_11978_ ( .A(\mreg/rf[11][5] ), .Z(\mreg/_04001_ ) );
BUF_X1 \mreg/_11979_ ( .A(\mreg/rf[10][5] ), .Z(\mreg/_03969_ ) );
BUF_X1 \mreg/_11980_ ( .A(\mreg/rf[9][5] ), .Z(\mreg/_04929_ ) );
BUF_X1 \mreg/_11981_ ( .A(\mreg/rf[8][5] ), .Z(\mreg/_04897_ ) );
BUF_X1 \mreg/_11982_ ( .A(\mreg/rf[7][5] ), .Z(\mreg/_04865_ ) );
BUF_X1 \mreg/_11983_ ( .A(\mreg/rf[6][5] ), .Z(\mreg/_04833_ ) );
BUF_X1 \mreg/_11984_ ( .A(\mreg/rf[5][5] ), .Z(\mreg/_04801_ ) );
BUF_X1 \mreg/_11985_ ( .A(\mreg/rf[4][5] ), .Z(\mreg/_04769_ ) );
BUF_X1 \mreg/_11986_ ( .A(\mreg/rf[3][5] ), .Z(\mreg/_04737_ ) );
BUF_X1 \mreg/_11987_ ( .A(\mreg/rf[2][5] ), .Z(\mreg/_04641_ ) );
BUF_X1 \mreg/_11988_ ( .A(\mreg/rf[1][5] ), .Z(\mreg/_04289_ ) );
BUF_X1 \mreg/_11989_ ( .A(\mreg/_03937_ ), .Z(\mem_wdata[5] ) );
BUF_X1 \mreg/_11990_ ( .A(\mreg/_00005_ ), .Z(\mreg/_00036_ ) );
BUF_X1 \mreg/_11991_ ( .A(\mreg/rf[30][6] ), .Z(\mreg/_04674_ ) );
BUF_X1 \mreg/_11992_ ( .A(\mreg/rf[29][6] ), .Z(\mreg/_04610_ ) );
BUF_X1 \mreg/_11993_ ( .A(\mreg/rf[28][6] ), .Z(\mreg/_04578_ ) );
BUF_X1 \mreg/_11994_ ( .A(\mreg/rf[27][6] ), .Z(\mreg/_04546_ ) );
BUF_X1 \mreg/_11995_ ( .A(\mreg/rf[26][6] ), .Z(\mreg/_04514_ ) );
BUF_X1 \mreg/_11996_ ( .A(\mreg/rf[25][6] ), .Z(\mreg/_04482_ ) );
BUF_X1 \mreg/_11997_ ( .A(\mreg/rf[24][6] ), .Z(\mreg/_04450_ ) );
BUF_X1 \mreg/_11998_ ( .A(\mreg/rf[23][6] ), .Z(\mreg/_04418_ ) );
BUF_X1 \mreg/_11999_ ( .A(\mreg/rf[22][6] ), .Z(\mreg/_04386_ ) );
BUF_X1 \mreg/_12000_ ( .A(\mreg/rf[21][6] ), .Z(\mreg/_04354_ ) );
BUF_X1 \mreg/_12001_ ( .A(\mreg/rf[20][6] ), .Z(\mreg/_04322_ ) );
BUF_X1 \mreg/_12002_ ( .A(\mreg/rf[19][6] ), .Z(\mreg/_04258_ ) );
BUF_X1 \mreg/_12003_ ( .A(\mreg/rf[18][6] ), .Z(\mreg/_04226_ ) );
BUF_X1 \mreg/_12004_ ( .A(\mreg/rf[17][6] ), .Z(\mreg/_04194_ ) );
BUF_X1 \mreg/_12005_ ( .A(\mreg/rf[16][6] ), .Z(\mreg/_04162_ ) );
BUF_X1 \mreg/_12006_ ( .A(\mreg/rf[15][6] ), .Z(\mreg/_04130_ ) );
BUF_X1 \mreg/_12007_ ( .A(\mreg/rf[14][6] ), .Z(\mreg/_04098_ ) );
BUF_X1 \mreg/_12008_ ( .A(\mreg/rf[13][6] ), .Z(\mreg/_04066_ ) );
BUF_X1 \mreg/_12009_ ( .A(\mreg/rf[12][6] ), .Z(\mreg/_04034_ ) );
BUF_X1 \mreg/_12010_ ( .A(\mreg/rf[11][6] ), .Z(\mreg/_04002_ ) );
BUF_X1 \mreg/_12011_ ( .A(\mreg/rf[10][6] ), .Z(\mreg/_03970_ ) );
BUF_X1 \mreg/_12012_ ( .A(\mreg/rf[9][6] ), .Z(\mreg/_04930_ ) );
BUF_X1 \mreg/_12013_ ( .A(\mreg/rf[8][6] ), .Z(\mreg/_04898_ ) );
BUF_X1 \mreg/_12014_ ( .A(\mreg/rf[7][6] ), .Z(\mreg/_04866_ ) );
BUF_X1 \mreg/_12015_ ( .A(\mreg/rf[6][6] ), .Z(\mreg/_04834_ ) );
BUF_X1 \mreg/_12016_ ( .A(\mreg/rf[5][6] ), .Z(\mreg/_04802_ ) );
BUF_X1 \mreg/_12017_ ( .A(\mreg/rf[4][6] ), .Z(\mreg/_04770_ ) );
BUF_X1 \mreg/_12018_ ( .A(\mreg/rf[3][6] ), .Z(\mreg/_04738_ ) );
BUF_X1 \mreg/_12019_ ( .A(\mreg/rf[2][6] ), .Z(\mreg/_04642_ ) );
BUF_X1 \mreg/_12020_ ( .A(\mreg/rf[1][6] ), .Z(\mreg/_04290_ ) );
BUF_X1 \mreg/_12021_ ( .A(\mreg/_03938_ ), .Z(\mem_wdata[6] ) );
BUF_X1 \mreg/_12022_ ( .A(\mreg/_00006_ ), .Z(\mreg/_00037_ ) );
BUF_X1 \mreg/_12023_ ( .A(\mreg/rf[30][7] ), .Z(\mreg/_04675_ ) );
BUF_X1 \mreg/_12024_ ( .A(\mreg/rf[29][7] ), .Z(\mreg/_04611_ ) );
BUF_X1 \mreg/_12025_ ( .A(\mreg/rf[28][7] ), .Z(\mreg/_04579_ ) );
BUF_X1 \mreg/_12026_ ( .A(\mreg/rf[27][7] ), .Z(\mreg/_04547_ ) );
BUF_X1 \mreg/_12027_ ( .A(\mreg/rf[26][7] ), .Z(\mreg/_04515_ ) );
BUF_X1 \mreg/_12028_ ( .A(\mreg/rf[25][7] ), .Z(\mreg/_04483_ ) );
BUF_X1 \mreg/_12029_ ( .A(\mreg/rf[24][7] ), .Z(\mreg/_04451_ ) );
BUF_X1 \mreg/_12030_ ( .A(\mreg/rf[23][7] ), .Z(\mreg/_04419_ ) );
BUF_X1 \mreg/_12031_ ( .A(\mreg/rf[22][7] ), .Z(\mreg/_04387_ ) );
BUF_X1 \mreg/_12032_ ( .A(\mreg/rf[21][7] ), .Z(\mreg/_04355_ ) );
BUF_X1 \mreg/_12033_ ( .A(\mreg/rf[20][7] ), .Z(\mreg/_04323_ ) );
BUF_X1 \mreg/_12034_ ( .A(\mreg/rf[19][7] ), .Z(\mreg/_04259_ ) );
BUF_X1 \mreg/_12035_ ( .A(\mreg/rf[18][7] ), .Z(\mreg/_04227_ ) );
BUF_X1 \mreg/_12036_ ( .A(\mreg/rf[17][7] ), .Z(\mreg/_04195_ ) );
BUF_X1 \mreg/_12037_ ( .A(\mreg/rf[16][7] ), .Z(\mreg/_04163_ ) );
BUF_X1 \mreg/_12038_ ( .A(\mreg/rf[15][7] ), .Z(\mreg/_04131_ ) );
BUF_X1 \mreg/_12039_ ( .A(\mreg/rf[14][7] ), .Z(\mreg/_04099_ ) );
BUF_X1 \mreg/_12040_ ( .A(\mreg/rf[13][7] ), .Z(\mreg/_04067_ ) );
BUF_X1 \mreg/_12041_ ( .A(\mreg/rf[12][7] ), .Z(\mreg/_04035_ ) );
BUF_X1 \mreg/_12042_ ( .A(\mreg/rf[11][7] ), .Z(\mreg/_04003_ ) );
BUF_X1 \mreg/_12043_ ( .A(\mreg/rf[10][7] ), .Z(\mreg/_03971_ ) );
BUF_X1 \mreg/_12044_ ( .A(\mreg/rf[9][7] ), .Z(\mreg/_04931_ ) );
BUF_X1 \mreg/_12045_ ( .A(\mreg/rf[8][7] ), .Z(\mreg/_04899_ ) );
BUF_X1 \mreg/_12046_ ( .A(\mreg/rf[7][7] ), .Z(\mreg/_04867_ ) );
BUF_X1 \mreg/_12047_ ( .A(\mreg/rf[6][7] ), .Z(\mreg/_04835_ ) );
BUF_X1 \mreg/_12048_ ( .A(\mreg/rf[5][7] ), .Z(\mreg/_04803_ ) );
BUF_X1 \mreg/_12049_ ( .A(\mreg/rf[4][7] ), .Z(\mreg/_04771_ ) );
BUF_X1 \mreg/_12050_ ( .A(\mreg/rf[3][7] ), .Z(\mreg/_04739_ ) );
BUF_X1 \mreg/_12051_ ( .A(\mreg/rf[2][7] ), .Z(\mreg/_04643_ ) );
BUF_X1 \mreg/_12052_ ( .A(\mreg/rf[1][7] ), .Z(\mreg/_04291_ ) );
BUF_X1 \mreg/_12053_ ( .A(\mreg/_03939_ ), .Z(\mem_wdata[7] ) );
BUF_X1 \mreg/_12054_ ( .A(\mreg/_00007_ ), .Z(\mreg/_00038_ ) );
BUF_X1 \mreg/_12055_ ( .A(\mreg/rf[30][8] ), .Z(\mreg/_04676_ ) );
BUF_X1 \mreg/_12056_ ( .A(\mreg/rf[29][8] ), .Z(\mreg/_04612_ ) );
BUF_X1 \mreg/_12057_ ( .A(\mreg/rf[28][8] ), .Z(\mreg/_04580_ ) );
BUF_X1 \mreg/_12058_ ( .A(\mreg/rf[27][8] ), .Z(\mreg/_04548_ ) );
BUF_X1 \mreg/_12059_ ( .A(\mreg/rf[26][8] ), .Z(\mreg/_04516_ ) );
BUF_X1 \mreg/_12060_ ( .A(\mreg/rf[25][8] ), .Z(\mreg/_04484_ ) );
BUF_X1 \mreg/_12061_ ( .A(\mreg/rf[24][8] ), .Z(\mreg/_04452_ ) );
BUF_X1 \mreg/_12062_ ( .A(\mreg/rf[23][8] ), .Z(\mreg/_04420_ ) );
BUF_X1 \mreg/_12063_ ( .A(\mreg/rf[22][8] ), .Z(\mreg/_04388_ ) );
BUF_X1 \mreg/_12064_ ( .A(\mreg/rf[21][8] ), .Z(\mreg/_04356_ ) );
BUF_X1 \mreg/_12065_ ( .A(\mreg/rf[20][8] ), .Z(\mreg/_04324_ ) );
BUF_X1 \mreg/_12066_ ( .A(\mreg/rf[19][8] ), .Z(\mreg/_04260_ ) );
BUF_X1 \mreg/_12067_ ( .A(\mreg/rf[18][8] ), .Z(\mreg/_04228_ ) );
BUF_X1 \mreg/_12068_ ( .A(\mreg/rf[17][8] ), .Z(\mreg/_04196_ ) );
BUF_X1 \mreg/_12069_ ( .A(\mreg/rf[16][8] ), .Z(\mreg/_04164_ ) );
BUF_X1 \mreg/_12070_ ( .A(\mreg/rf[15][8] ), .Z(\mreg/_04132_ ) );
BUF_X1 \mreg/_12071_ ( .A(\mreg/rf[14][8] ), .Z(\mreg/_04100_ ) );
BUF_X1 \mreg/_12072_ ( .A(\mreg/rf[13][8] ), .Z(\mreg/_04068_ ) );
BUF_X1 \mreg/_12073_ ( .A(\mreg/rf[12][8] ), .Z(\mreg/_04036_ ) );
BUF_X1 \mreg/_12074_ ( .A(\mreg/rf[11][8] ), .Z(\mreg/_04004_ ) );
BUF_X1 \mreg/_12075_ ( .A(\mreg/rf[10][8] ), .Z(\mreg/_03972_ ) );
BUF_X1 \mreg/_12076_ ( .A(\mreg/rf[9][8] ), .Z(\mreg/_04932_ ) );
BUF_X1 \mreg/_12077_ ( .A(\mreg/rf[8][8] ), .Z(\mreg/_04900_ ) );
BUF_X1 \mreg/_12078_ ( .A(\mreg/rf[7][8] ), .Z(\mreg/_04868_ ) );
BUF_X1 \mreg/_12079_ ( .A(\mreg/rf[6][8] ), .Z(\mreg/_04836_ ) );
BUF_X1 \mreg/_12080_ ( .A(\mreg/rf[5][8] ), .Z(\mreg/_04804_ ) );
BUF_X1 \mreg/_12081_ ( .A(\mreg/rf[4][8] ), .Z(\mreg/_04772_ ) );
BUF_X1 \mreg/_12082_ ( .A(\mreg/rf[3][8] ), .Z(\mreg/_04740_ ) );
BUF_X1 \mreg/_12083_ ( .A(\mreg/rf[2][8] ), .Z(\mreg/_04644_ ) );
BUF_X1 \mreg/_12084_ ( .A(\mreg/rf[1][8] ), .Z(\mreg/_04292_ ) );
BUF_X1 \mreg/_12085_ ( .A(\mreg/_03940_ ), .Z(\mem_wdata[8] ) );
BUF_X1 \mreg/_12086_ ( .A(\mreg/_00008_ ), .Z(\mreg/_00039_ ) );
BUF_X1 \mreg/_12087_ ( .A(\mreg/rf[30][9] ), .Z(\mreg/_04677_ ) );
BUF_X1 \mreg/_12088_ ( .A(\mreg/rf[29][9] ), .Z(\mreg/_04613_ ) );
BUF_X1 \mreg/_12089_ ( .A(\mreg/rf[28][9] ), .Z(\mreg/_04581_ ) );
BUF_X1 \mreg/_12090_ ( .A(\mreg/rf[27][9] ), .Z(\mreg/_04549_ ) );
BUF_X1 \mreg/_12091_ ( .A(\mreg/rf[26][9] ), .Z(\mreg/_04517_ ) );
BUF_X1 \mreg/_12092_ ( .A(\mreg/rf[25][9] ), .Z(\mreg/_04485_ ) );
BUF_X1 \mreg/_12093_ ( .A(\mreg/rf[24][9] ), .Z(\mreg/_04453_ ) );
BUF_X1 \mreg/_12094_ ( .A(\mreg/rf[23][9] ), .Z(\mreg/_04421_ ) );
BUF_X1 \mreg/_12095_ ( .A(\mreg/rf[22][9] ), .Z(\mreg/_04389_ ) );
BUF_X1 \mreg/_12096_ ( .A(\mreg/rf[21][9] ), .Z(\mreg/_04357_ ) );
BUF_X1 \mreg/_12097_ ( .A(\mreg/rf[20][9] ), .Z(\mreg/_04325_ ) );
BUF_X1 \mreg/_12098_ ( .A(\mreg/rf[19][9] ), .Z(\mreg/_04261_ ) );
BUF_X1 \mreg/_12099_ ( .A(\mreg/rf[18][9] ), .Z(\mreg/_04229_ ) );
BUF_X1 \mreg/_12100_ ( .A(\mreg/rf[17][9] ), .Z(\mreg/_04197_ ) );
BUF_X1 \mreg/_12101_ ( .A(\mreg/rf[16][9] ), .Z(\mreg/_04165_ ) );
BUF_X1 \mreg/_12102_ ( .A(\mreg/rf[15][9] ), .Z(\mreg/_04133_ ) );
BUF_X1 \mreg/_12103_ ( .A(\mreg/rf[14][9] ), .Z(\mreg/_04101_ ) );
BUF_X1 \mreg/_12104_ ( .A(\mreg/rf[13][9] ), .Z(\mreg/_04069_ ) );
BUF_X1 \mreg/_12105_ ( .A(\mreg/rf[12][9] ), .Z(\mreg/_04037_ ) );
BUF_X1 \mreg/_12106_ ( .A(\mreg/rf[11][9] ), .Z(\mreg/_04005_ ) );
BUF_X1 \mreg/_12107_ ( .A(\mreg/rf[10][9] ), .Z(\mreg/_03973_ ) );
BUF_X1 \mreg/_12108_ ( .A(\mreg/rf[9][9] ), .Z(\mreg/_04933_ ) );
BUF_X1 \mreg/_12109_ ( .A(\mreg/rf[8][9] ), .Z(\mreg/_04901_ ) );
BUF_X1 \mreg/_12110_ ( .A(\mreg/rf[7][9] ), .Z(\mreg/_04869_ ) );
BUF_X1 \mreg/_12111_ ( .A(\mreg/rf[6][9] ), .Z(\mreg/_04837_ ) );
BUF_X1 \mreg/_12112_ ( .A(\mreg/rf[5][9] ), .Z(\mreg/_04805_ ) );
BUF_X1 \mreg/_12113_ ( .A(\mreg/rf[4][9] ), .Z(\mreg/_04773_ ) );
BUF_X1 \mreg/_12114_ ( .A(\mreg/rf[3][9] ), .Z(\mreg/_04741_ ) );
BUF_X1 \mreg/_12115_ ( .A(\mreg/rf[2][9] ), .Z(\mreg/_04645_ ) );
BUF_X1 \mreg/_12116_ ( .A(\mreg/rf[1][9] ), .Z(\mreg/_04293_ ) );
BUF_X1 \mreg/_12117_ ( .A(\mreg/_03941_ ), .Z(\mem_wdata[9] ) );
BUF_X1 \mreg/_12118_ ( .A(\mreg/_00009_ ), .Z(\mreg/_00040_ ) );
BUF_X1 \mreg/_12119_ ( .A(\mreg/rf[30][10] ), .Z(\mreg/_04647_ ) );
BUF_X1 \mreg/_12120_ ( .A(\mreg/rf[29][10] ), .Z(\mreg/_04583_ ) );
BUF_X1 \mreg/_12121_ ( .A(\mreg/rf[28][10] ), .Z(\mreg/_04551_ ) );
BUF_X1 \mreg/_12122_ ( .A(\mreg/rf[27][10] ), .Z(\mreg/_04519_ ) );
BUF_X1 \mreg/_12123_ ( .A(\mreg/rf[26][10] ), .Z(\mreg/_04487_ ) );
BUF_X1 \mreg/_12124_ ( .A(\mreg/rf[25][10] ), .Z(\mreg/_04455_ ) );
BUF_X1 \mreg/_12125_ ( .A(\mreg/rf[24][10] ), .Z(\mreg/_04423_ ) );
BUF_X1 \mreg/_12126_ ( .A(\mreg/rf[23][10] ), .Z(\mreg/_04391_ ) );
BUF_X1 \mreg/_12127_ ( .A(\mreg/rf[22][10] ), .Z(\mreg/_04359_ ) );
BUF_X1 \mreg/_12128_ ( .A(\mreg/rf[21][10] ), .Z(\mreg/_04327_ ) );
BUF_X1 \mreg/_12129_ ( .A(\mreg/rf[20][10] ), .Z(\mreg/_04295_ ) );
BUF_X1 \mreg/_12130_ ( .A(\mreg/rf[19][10] ), .Z(\mreg/_04231_ ) );
BUF_X1 \mreg/_12131_ ( .A(\mreg/rf[18][10] ), .Z(\mreg/_04199_ ) );
BUF_X1 \mreg/_12132_ ( .A(\mreg/rf[17][10] ), .Z(\mreg/_04167_ ) );
BUF_X1 \mreg/_12133_ ( .A(\mreg/rf[16][10] ), .Z(\mreg/_04135_ ) );
BUF_X1 \mreg/_12134_ ( .A(\mreg/rf[15][10] ), .Z(\mreg/_04103_ ) );
BUF_X1 \mreg/_12135_ ( .A(\mreg/rf[14][10] ), .Z(\mreg/_04071_ ) );
BUF_X1 \mreg/_12136_ ( .A(\mreg/rf[13][10] ), .Z(\mreg/_04039_ ) );
BUF_X1 \mreg/_12137_ ( .A(\mreg/rf[12][10] ), .Z(\mreg/_04007_ ) );
BUF_X1 \mreg/_12138_ ( .A(\mreg/rf[11][10] ), .Z(\mreg/_03975_ ) );
BUF_X1 \mreg/_12139_ ( .A(\mreg/rf[10][10] ), .Z(\mreg/_03943_ ) );
BUF_X1 \mreg/_12140_ ( .A(\mreg/rf[9][10] ), .Z(\mreg/_04903_ ) );
BUF_X1 \mreg/_12141_ ( .A(\mreg/rf[8][10] ), .Z(\mreg/_04871_ ) );
BUF_X1 \mreg/_12142_ ( .A(\mreg/rf[7][10] ), .Z(\mreg/_04839_ ) );
BUF_X1 \mreg/_12143_ ( .A(\mreg/rf[6][10] ), .Z(\mreg/_04807_ ) );
BUF_X1 \mreg/_12144_ ( .A(\mreg/rf[5][10] ), .Z(\mreg/_04775_ ) );
BUF_X1 \mreg/_12145_ ( .A(\mreg/rf[4][10] ), .Z(\mreg/_04743_ ) );
BUF_X1 \mreg/_12146_ ( .A(\mreg/rf[3][10] ), .Z(\mreg/_04711_ ) );
BUF_X1 \mreg/_12147_ ( .A(\mreg/rf[2][10] ), .Z(\mreg/_04615_ ) );
BUF_X1 \mreg/_12148_ ( .A(\mreg/rf[1][10] ), .Z(\mreg/_04263_ ) );
BUF_X1 \mreg/_12149_ ( .A(\mreg/_03911_ ), .Z(\mem_wdata[10] ) );
BUF_X1 \mreg/_12150_ ( .A(\mreg/_00010_ ), .Z(\mreg/_00041_ ) );
BUF_X1 \mreg/_12151_ ( .A(\mreg/rf[30][11] ), .Z(\mreg/_04648_ ) );
BUF_X1 \mreg/_12152_ ( .A(\mreg/rf[29][11] ), .Z(\mreg/_04584_ ) );
BUF_X1 \mreg/_12153_ ( .A(\mreg/rf[28][11] ), .Z(\mreg/_04552_ ) );
BUF_X1 \mreg/_12154_ ( .A(\mreg/rf[27][11] ), .Z(\mreg/_04520_ ) );
BUF_X1 \mreg/_12155_ ( .A(\mreg/rf[26][11] ), .Z(\mreg/_04488_ ) );
BUF_X1 \mreg/_12156_ ( .A(\mreg/rf[25][11] ), .Z(\mreg/_04456_ ) );
BUF_X1 \mreg/_12157_ ( .A(\mreg/rf[24][11] ), .Z(\mreg/_04424_ ) );
BUF_X1 \mreg/_12158_ ( .A(\mreg/rf[23][11] ), .Z(\mreg/_04392_ ) );
BUF_X1 \mreg/_12159_ ( .A(\mreg/rf[22][11] ), .Z(\mreg/_04360_ ) );
BUF_X1 \mreg/_12160_ ( .A(\mreg/rf[21][11] ), .Z(\mreg/_04328_ ) );
BUF_X1 \mreg/_12161_ ( .A(\mreg/rf[20][11] ), .Z(\mreg/_04296_ ) );
BUF_X1 \mreg/_12162_ ( .A(\mreg/rf[19][11] ), .Z(\mreg/_04232_ ) );
BUF_X1 \mreg/_12163_ ( .A(\mreg/rf[18][11] ), .Z(\mreg/_04200_ ) );
BUF_X1 \mreg/_12164_ ( .A(\mreg/rf[17][11] ), .Z(\mreg/_04168_ ) );
BUF_X1 \mreg/_12165_ ( .A(\mreg/rf[16][11] ), .Z(\mreg/_04136_ ) );
BUF_X1 \mreg/_12166_ ( .A(\mreg/rf[15][11] ), .Z(\mreg/_04104_ ) );
BUF_X1 \mreg/_12167_ ( .A(\mreg/rf[14][11] ), .Z(\mreg/_04072_ ) );
BUF_X1 \mreg/_12168_ ( .A(\mreg/rf[13][11] ), .Z(\mreg/_04040_ ) );
BUF_X1 \mreg/_12169_ ( .A(\mreg/rf[12][11] ), .Z(\mreg/_04008_ ) );
BUF_X1 \mreg/_12170_ ( .A(\mreg/rf[11][11] ), .Z(\mreg/_03976_ ) );
BUF_X1 \mreg/_12171_ ( .A(\mreg/rf[10][11] ), .Z(\mreg/_03944_ ) );
BUF_X1 \mreg/_12172_ ( .A(\mreg/rf[9][11] ), .Z(\mreg/_04904_ ) );
BUF_X1 \mreg/_12173_ ( .A(\mreg/rf[8][11] ), .Z(\mreg/_04872_ ) );
BUF_X1 \mreg/_12174_ ( .A(\mreg/rf[7][11] ), .Z(\mreg/_04840_ ) );
BUF_X1 \mreg/_12175_ ( .A(\mreg/rf[6][11] ), .Z(\mreg/_04808_ ) );
BUF_X1 \mreg/_12176_ ( .A(\mreg/rf[5][11] ), .Z(\mreg/_04776_ ) );
BUF_X1 \mreg/_12177_ ( .A(\mreg/rf[4][11] ), .Z(\mreg/_04744_ ) );
BUF_X1 \mreg/_12178_ ( .A(\mreg/rf[3][11] ), .Z(\mreg/_04712_ ) );
BUF_X1 \mreg/_12179_ ( .A(\mreg/rf[2][11] ), .Z(\mreg/_04616_ ) );
BUF_X1 \mreg/_12180_ ( .A(\mreg/rf[1][11] ), .Z(\mreg/_04264_ ) );
BUF_X1 \mreg/_12181_ ( .A(\mreg/_03912_ ), .Z(\mem_wdata[11] ) );
BUF_X1 \mreg/_12182_ ( .A(\mreg/_00011_ ), .Z(\mreg/_00042_ ) );
BUF_X1 \mreg/_12183_ ( .A(\mreg/rf[30][12] ), .Z(\mreg/_04649_ ) );
BUF_X1 \mreg/_12184_ ( .A(\mreg/rf[29][12] ), .Z(\mreg/_04585_ ) );
BUF_X1 \mreg/_12185_ ( .A(\mreg/rf[28][12] ), .Z(\mreg/_04553_ ) );
BUF_X1 \mreg/_12186_ ( .A(\mreg/rf[27][12] ), .Z(\mreg/_04521_ ) );
BUF_X1 \mreg/_12187_ ( .A(\mreg/rf[26][12] ), .Z(\mreg/_04489_ ) );
BUF_X1 \mreg/_12188_ ( .A(\mreg/rf[25][12] ), .Z(\mreg/_04457_ ) );
BUF_X1 \mreg/_12189_ ( .A(\mreg/rf[24][12] ), .Z(\mreg/_04425_ ) );
BUF_X1 \mreg/_12190_ ( .A(\mreg/rf[23][12] ), .Z(\mreg/_04393_ ) );
BUF_X1 \mreg/_12191_ ( .A(\mreg/rf[22][12] ), .Z(\mreg/_04361_ ) );
BUF_X1 \mreg/_12192_ ( .A(\mreg/rf[21][12] ), .Z(\mreg/_04329_ ) );
BUF_X1 \mreg/_12193_ ( .A(\mreg/rf[20][12] ), .Z(\mreg/_04297_ ) );
BUF_X1 \mreg/_12194_ ( .A(\mreg/rf[19][12] ), .Z(\mreg/_04233_ ) );
BUF_X1 \mreg/_12195_ ( .A(\mreg/rf[18][12] ), .Z(\mreg/_04201_ ) );
BUF_X1 \mreg/_12196_ ( .A(\mreg/rf[17][12] ), .Z(\mreg/_04169_ ) );
BUF_X1 \mreg/_12197_ ( .A(\mreg/rf[16][12] ), .Z(\mreg/_04137_ ) );
BUF_X1 \mreg/_12198_ ( .A(\mreg/rf[15][12] ), .Z(\mreg/_04105_ ) );
BUF_X1 \mreg/_12199_ ( .A(\mreg/rf[14][12] ), .Z(\mreg/_04073_ ) );
BUF_X1 \mreg/_12200_ ( .A(\mreg/rf[13][12] ), .Z(\mreg/_04041_ ) );
BUF_X1 \mreg/_12201_ ( .A(\mreg/rf[12][12] ), .Z(\mreg/_04009_ ) );
BUF_X1 \mreg/_12202_ ( .A(\mreg/rf[11][12] ), .Z(\mreg/_03977_ ) );
BUF_X1 \mreg/_12203_ ( .A(\mreg/rf[10][12] ), .Z(\mreg/_03945_ ) );
BUF_X1 \mreg/_12204_ ( .A(\mreg/rf[9][12] ), .Z(\mreg/_04905_ ) );
BUF_X1 \mreg/_12205_ ( .A(\mreg/rf[8][12] ), .Z(\mreg/_04873_ ) );
BUF_X1 \mreg/_12206_ ( .A(\mreg/rf[7][12] ), .Z(\mreg/_04841_ ) );
BUF_X1 \mreg/_12207_ ( .A(\mreg/rf[6][12] ), .Z(\mreg/_04809_ ) );
BUF_X1 \mreg/_12208_ ( .A(\mreg/rf[5][12] ), .Z(\mreg/_04777_ ) );
BUF_X1 \mreg/_12209_ ( .A(\mreg/rf[4][12] ), .Z(\mreg/_04745_ ) );
BUF_X1 \mreg/_12210_ ( .A(\mreg/rf[3][12] ), .Z(\mreg/_04713_ ) );
BUF_X1 \mreg/_12211_ ( .A(\mreg/rf[2][12] ), .Z(\mreg/_04617_ ) );
BUF_X1 \mreg/_12212_ ( .A(\mreg/rf[1][12] ), .Z(\mreg/_04265_ ) );
BUF_X1 \mreg/_12213_ ( .A(\mreg/_03913_ ), .Z(\mem_wdata[12] ) );
BUF_X1 \mreg/_12214_ ( .A(\mreg/_00012_ ), .Z(\mreg/_00043_ ) );
BUF_X1 \mreg/_12215_ ( .A(\mreg/rf[30][13] ), .Z(\mreg/_04650_ ) );
BUF_X1 \mreg/_12216_ ( .A(\mreg/rf[29][13] ), .Z(\mreg/_04586_ ) );
BUF_X1 \mreg/_12217_ ( .A(\mreg/rf[28][13] ), .Z(\mreg/_04554_ ) );
BUF_X1 \mreg/_12218_ ( .A(\mreg/rf[27][13] ), .Z(\mreg/_04522_ ) );
BUF_X1 \mreg/_12219_ ( .A(\mreg/rf[26][13] ), .Z(\mreg/_04490_ ) );
BUF_X1 \mreg/_12220_ ( .A(\mreg/rf[25][13] ), .Z(\mreg/_04458_ ) );
BUF_X1 \mreg/_12221_ ( .A(\mreg/rf[24][13] ), .Z(\mreg/_04426_ ) );
BUF_X1 \mreg/_12222_ ( .A(\mreg/rf[23][13] ), .Z(\mreg/_04394_ ) );
BUF_X1 \mreg/_12223_ ( .A(\mreg/rf[22][13] ), .Z(\mreg/_04362_ ) );
BUF_X1 \mreg/_12224_ ( .A(\mreg/rf[21][13] ), .Z(\mreg/_04330_ ) );
BUF_X1 \mreg/_12225_ ( .A(\mreg/rf[20][13] ), .Z(\mreg/_04298_ ) );
BUF_X1 \mreg/_12226_ ( .A(\mreg/rf[19][13] ), .Z(\mreg/_04234_ ) );
BUF_X1 \mreg/_12227_ ( .A(\mreg/rf[18][13] ), .Z(\mreg/_04202_ ) );
BUF_X1 \mreg/_12228_ ( .A(\mreg/rf[17][13] ), .Z(\mreg/_04170_ ) );
BUF_X1 \mreg/_12229_ ( .A(\mreg/rf[16][13] ), .Z(\mreg/_04138_ ) );
BUF_X1 \mreg/_12230_ ( .A(\mreg/rf[15][13] ), .Z(\mreg/_04106_ ) );
BUF_X1 \mreg/_12231_ ( .A(\mreg/rf[14][13] ), .Z(\mreg/_04074_ ) );
BUF_X1 \mreg/_12232_ ( .A(\mreg/rf[13][13] ), .Z(\mreg/_04042_ ) );
BUF_X1 \mreg/_12233_ ( .A(\mreg/rf[12][13] ), .Z(\mreg/_04010_ ) );
BUF_X1 \mreg/_12234_ ( .A(\mreg/rf[11][13] ), .Z(\mreg/_03978_ ) );
BUF_X1 \mreg/_12235_ ( .A(\mreg/rf[10][13] ), .Z(\mreg/_03946_ ) );
BUF_X1 \mreg/_12236_ ( .A(\mreg/rf[9][13] ), .Z(\mreg/_04906_ ) );
BUF_X1 \mreg/_12237_ ( .A(\mreg/rf[8][13] ), .Z(\mreg/_04874_ ) );
BUF_X1 \mreg/_12238_ ( .A(\mreg/rf[7][13] ), .Z(\mreg/_04842_ ) );
BUF_X1 \mreg/_12239_ ( .A(\mreg/rf[6][13] ), .Z(\mreg/_04810_ ) );
BUF_X1 \mreg/_12240_ ( .A(\mreg/rf[5][13] ), .Z(\mreg/_04778_ ) );
BUF_X1 \mreg/_12241_ ( .A(\mreg/rf[4][13] ), .Z(\mreg/_04746_ ) );
BUF_X1 \mreg/_12242_ ( .A(\mreg/rf[3][13] ), .Z(\mreg/_04714_ ) );
BUF_X1 \mreg/_12243_ ( .A(\mreg/rf[2][13] ), .Z(\mreg/_04618_ ) );
BUF_X1 \mreg/_12244_ ( .A(\mreg/rf[1][13] ), .Z(\mreg/_04266_ ) );
BUF_X1 \mreg/_12245_ ( .A(\mreg/_03914_ ), .Z(\mem_wdata[13] ) );
BUF_X1 \mreg/_12246_ ( .A(\mreg/_00013_ ), .Z(\mreg/_00044_ ) );
BUF_X1 \mreg/_12247_ ( .A(\mreg/rf[30][14] ), .Z(\mreg/_04651_ ) );
BUF_X1 \mreg/_12248_ ( .A(\mreg/rf[29][14] ), .Z(\mreg/_04587_ ) );
BUF_X1 \mreg/_12249_ ( .A(\mreg/rf[28][14] ), .Z(\mreg/_04555_ ) );
BUF_X1 \mreg/_12250_ ( .A(\mreg/rf[27][14] ), .Z(\mreg/_04523_ ) );
BUF_X1 \mreg/_12251_ ( .A(\mreg/rf[26][14] ), .Z(\mreg/_04491_ ) );
BUF_X1 \mreg/_12252_ ( .A(\mreg/rf[25][14] ), .Z(\mreg/_04459_ ) );
BUF_X1 \mreg/_12253_ ( .A(\mreg/rf[24][14] ), .Z(\mreg/_04427_ ) );
BUF_X1 \mreg/_12254_ ( .A(\mreg/rf[23][14] ), .Z(\mreg/_04395_ ) );
BUF_X1 \mreg/_12255_ ( .A(\mreg/rf[22][14] ), .Z(\mreg/_04363_ ) );
BUF_X1 \mreg/_12256_ ( .A(\mreg/rf[21][14] ), .Z(\mreg/_04331_ ) );
BUF_X1 \mreg/_12257_ ( .A(\mreg/rf[20][14] ), .Z(\mreg/_04299_ ) );
BUF_X1 \mreg/_12258_ ( .A(\mreg/rf[19][14] ), .Z(\mreg/_04235_ ) );
BUF_X1 \mreg/_12259_ ( .A(\mreg/rf[18][14] ), .Z(\mreg/_04203_ ) );
BUF_X1 \mreg/_12260_ ( .A(\mreg/rf[17][14] ), .Z(\mreg/_04171_ ) );
BUF_X1 \mreg/_12261_ ( .A(\mreg/rf[16][14] ), .Z(\mreg/_04139_ ) );
BUF_X1 \mreg/_12262_ ( .A(\mreg/rf[15][14] ), .Z(\mreg/_04107_ ) );
BUF_X1 \mreg/_12263_ ( .A(\mreg/rf[14][14] ), .Z(\mreg/_04075_ ) );
BUF_X1 \mreg/_12264_ ( .A(\mreg/rf[13][14] ), .Z(\mreg/_04043_ ) );
BUF_X1 \mreg/_12265_ ( .A(\mreg/rf[12][14] ), .Z(\mreg/_04011_ ) );
BUF_X1 \mreg/_12266_ ( .A(\mreg/rf[11][14] ), .Z(\mreg/_03979_ ) );
BUF_X1 \mreg/_12267_ ( .A(\mreg/rf[10][14] ), .Z(\mreg/_03947_ ) );
BUF_X1 \mreg/_12268_ ( .A(\mreg/rf[9][14] ), .Z(\mreg/_04907_ ) );
BUF_X1 \mreg/_12269_ ( .A(\mreg/rf[8][14] ), .Z(\mreg/_04875_ ) );
BUF_X1 \mreg/_12270_ ( .A(\mreg/rf[7][14] ), .Z(\mreg/_04843_ ) );
BUF_X1 \mreg/_12271_ ( .A(\mreg/rf[6][14] ), .Z(\mreg/_04811_ ) );
BUF_X1 \mreg/_12272_ ( .A(\mreg/rf[5][14] ), .Z(\mreg/_04779_ ) );
BUF_X1 \mreg/_12273_ ( .A(\mreg/rf[4][14] ), .Z(\mreg/_04747_ ) );
BUF_X1 \mreg/_12274_ ( .A(\mreg/rf[3][14] ), .Z(\mreg/_04715_ ) );
BUF_X1 \mreg/_12275_ ( .A(\mreg/rf[2][14] ), .Z(\mreg/_04619_ ) );
BUF_X1 \mreg/_12276_ ( .A(\mreg/rf[1][14] ), .Z(\mreg/_04267_ ) );
BUF_X1 \mreg/_12277_ ( .A(\mreg/_03915_ ), .Z(\mem_wdata[14] ) );
BUF_X1 \mreg/_12278_ ( .A(\mreg/_00014_ ), .Z(\mreg/_00045_ ) );
BUF_X1 \mreg/_12279_ ( .A(\mreg/rf[30][15] ), .Z(\mreg/_04652_ ) );
BUF_X1 \mreg/_12280_ ( .A(\mreg/rf[29][15] ), .Z(\mreg/_04588_ ) );
BUF_X1 \mreg/_12281_ ( .A(\mreg/rf[28][15] ), .Z(\mreg/_04556_ ) );
BUF_X1 \mreg/_12282_ ( .A(\mreg/rf[27][15] ), .Z(\mreg/_04524_ ) );
BUF_X1 \mreg/_12283_ ( .A(\mreg/rf[26][15] ), .Z(\mreg/_04492_ ) );
BUF_X1 \mreg/_12284_ ( .A(\mreg/rf[25][15] ), .Z(\mreg/_04460_ ) );
BUF_X1 \mreg/_12285_ ( .A(\mreg/rf[24][15] ), .Z(\mreg/_04428_ ) );
BUF_X1 \mreg/_12286_ ( .A(\mreg/rf[23][15] ), .Z(\mreg/_04396_ ) );
BUF_X1 \mreg/_12287_ ( .A(\mreg/rf[22][15] ), .Z(\mreg/_04364_ ) );
BUF_X1 \mreg/_12288_ ( .A(\mreg/rf[21][15] ), .Z(\mreg/_04332_ ) );
BUF_X1 \mreg/_12289_ ( .A(\mreg/rf[20][15] ), .Z(\mreg/_04300_ ) );
BUF_X1 \mreg/_12290_ ( .A(\mreg/rf[19][15] ), .Z(\mreg/_04236_ ) );
BUF_X1 \mreg/_12291_ ( .A(\mreg/rf[18][15] ), .Z(\mreg/_04204_ ) );
BUF_X1 \mreg/_12292_ ( .A(\mreg/rf[17][15] ), .Z(\mreg/_04172_ ) );
BUF_X1 \mreg/_12293_ ( .A(\mreg/rf[16][15] ), .Z(\mreg/_04140_ ) );
BUF_X1 \mreg/_12294_ ( .A(\mreg/rf[15][15] ), .Z(\mreg/_04108_ ) );
BUF_X1 \mreg/_12295_ ( .A(\mreg/rf[14][15] ), .Z(\mreg/_04076_ ) );
BUF_X1 \mreg/_12296_ ( .A(\mreg/rf[13][15] ), .Z(\mreg/_04044_ ) );
BUF_X1 \mreg/_12297_ ( .A(\mreg/rf[12][15] ), .Z(\mreg/_04012_ ) );
BUF_X1 \mreg/_12298_ ( .A(\mreg/rf[11][15] ), .Z(\mreg/_03980_ ) );
BUF_X1 \mreg/_12299_ ( .A(\mreg/rf[10][15] ), .Z(\mreg/_03948_ ) );
BUF_X1 \mreg/_12300_ ( .A(\mreg/rf[9][15] ), .Z(\mreg/_04908_ ) );
BUF_X1 \mreg/_12301_ ( .A(\mreg/rf[8][15] ), .Z(\mreg/_04876_ ) );
BUF_X1 \mreg/_12302_ ( .A(\mreg/rf[7][15] ), .Z(\mreg/_04844_ ) );
BUF_X1 \mreg/_12303_ ( .A(\mreg/rf[6][15] ), .Z(\mreg/_04812_ ) );
BUF_X1 \mreg/_12304_ ( .A(\mreg/rf[5][15] ), .Z(\mreg/_04780_ ) );
BUF_X1 \mreg/_12305_ ( .A(\mreg/rf[4][15] ), .Z(\mreg/_04748_ ) );
BUF_X1 \mreg/_12306_ ( .A(\mreg/rf[3][15] ), .Z(\mreg/_04716_ ) );
BUF_X1 \mreg/_12307_ ( .A(\mreg/rf[2][15] ), .Z(\mreg/_04620_ ) );
BUF_X1 \mreg/_12308_ ( .A(\mreg/rf[1][15] ), .Z(\mreg/_04268_ ) );
BUF_X1 \mreg/_12309_ ( .A(\mreg/_03916_ ), .Z(\mem_wdata[15] ) );
BUF_X1 \mreg/_12310_ ( .A(\mreg/_00015_ ), .Z(\mreg/_00046_ ) );
BUF_X1 \mreg/_12311_ ( .A(\mreg/rf[30][16] ), .Z(\mreg/_04653_ ) );
BUF_X1 \mreg/_12312_ ( .A(\mreg/rf[29][16] ), .Z(\mreg/_04589_ ) );
BUF_X1 \mreg/_12313_ ( .A(\mreg/rf[28][16] ), .Z(\mreg/_04557_ ) );
BUF_X1 \mreg/_12314_ ( .A(\mreg/rf[27][16] ), .Z(\mreg/_04525_ ) );
BUF_X1 \mreg/_12315_ ( .A(\mreg/rf[26][16] ), .Z(\mreg/_04493_ ) );
BUF_X1 \mreg/_12316_ ( .A(\mreg/rf[25][16] ), .Z(\mreg/_04461_ ) );
BUF_X1 \mreg/_12317_ ( .A(\mreg/rf[24][16] ), .Z(\mreg/_04429_ ) );
BUF_X1 \mreg/_12318_ ( .A(\mreg/rf[23][16] ), .Z(\mreg/_04397_ ) );
BUF_X1 \mreg/_12319_ ( .A(\mreg/rf[22][16] ), .Z(\mreg/_04365_ ) );
BUF_X1 \mreg/_12320_ ( .A(\mreg/rf[21][16] ), .Z(\mreg/_04333_ ) );
BUF_X1 \mreg/_12321_ ( .A(\mreg/rf[20][16] ), .Z(\mreg/_04301_ ) );
BUF_X1 \mreg/_12322_ ( .A(\mreg/rf[19][16] ), .Z(\mreg/_04237_ ) );
BUF_X1 \mreg/_12323_ ( .A(\mreg/rf[18][16] ), .Z(\mreg/_04205_ ) );
BUF_X1 \mreg/_12324_ ( .A(\mreg/rf[17][16] ), .Z(\mreg/_04173_ ) );
BUF_X1 \mreg/_12325_ ( .A(\mreg/rf[16][16] ), .Z(\mreg/_04141_ ) );
BUF_X1 \mreg/_12326_ ( .A(\mreg/rf[15][16] ), .Z(\mreg/_04109_ ) );
BUF_X1 \mreg/_12327_ ( .A(\mreg/rf[14][16] ), .Z(\mreg/_04077_ ) );
BUF_X1 \mreg/_12328_ ( .A(\mreg/rf[13][16] ), .Z(\mreg/_04045_ ) );
BUF_X1 \mreg/_12329_ ( .A(\mreg/rf[12][16] ), .Z(\mreg/_04013_ ) );
BUF_X1 \mreg/_12330_ ( .A(\mreg/rf[11][16] ), .Z(\mreg/_03981_ ) );
BUF_X1 \mreg/_12331_ ( .A(\mreg/rf[10][16] ), .Z(\mreg/_03949_ ) );
BUF_X1 \mreg/_12332_ ( .A(\mreg/rf[9][16] ), .Z(\mreg/_04909_ ) );
BUF_X1 \mreg/_12333_ ( .A(\mreg/rf[8][16] ), .Z(\mreg/_04877_ ) );
BUF_X1 \mreg/_12334_ ( .A(\mreg/rf[7][16] ), .Z(\mreg/_04845_ ) );
BUF_X1 \mreg/_12335_ ( .A(\mreg/rf[6][16] ), .Z(\mreg/_04813_ ) );
BUF_X1 \mreg/_12336_ ( .A(\mreg/rf[5][16] ), .Z(\mreg/_04781_ ) );
BUF_X1 \mreg/_12337_ ( .A(\mreg/rf[4][16] ), .Z(\mreg/_04749_ ) );
BUF_X1 \mreg/_12338_ ( .A(\mreg/rf[3][16] ), .Z(\mreg/_04717_ ) );
BUF_X1 \mreg/_12339_ ( .A(\mreg/rf[2][16] ), .Z(\mreg/_04621_ ) );
BUF_X1 \mreg/_12340_ ( .A(\mreg/rf[1][16] ), .Z(\mreg/_04269_ ) );
BUF_X1 \mreg/_12341_ ( .A(\mreg/_03917_ ), .Z(\mem_wdata[16] ) );
BUF_X1 \mreg/_12342_ ( .A(\mreg/_00016_ ), .Z(\mreg/_00047_ ) );
BUF_X1 \mreg/_12343_ ( .A(\mreg/rf[30][17] ), .Z(\mreg/_04654_ ) );
BUF_X1 \mreg/_12344_ ( .A(\mreg/rf[29][17] ), .Z(\mreg/_04590_ ) );
BUF_X1 \mreg/_12345_ ( .A(\mreg/rf[28][17] ), .Z(\mreg/_04558_ ) );
BUF_X1 \mreg/_12346_ ( .A(\mreg/rf[27][17] ), .Z(\mreg/_04526_ ) );
BUF_X1 \mreg/_12347_ ( .A(\mreg/rf[26][17] ), .Z(\mreg/_04494_ ) );
BUF_X1 \mreg/_12348_ ( .A(\mreg/rf[25][17] ), .Z(\mreg/_04462_ ) );
BUF_X1 \mreg/_12349_ ( .A(\mreg/rf[24][17] ), .Z(\mreg/_04430_ ) );
BUF_X1 \mreg/_12350_ ( .A(\mreg/rf[23][17] ), .Z(\mreg/_04398_ ) );
BUF_X1 \mreg/_12351_ ( .A(\mreg/rf[22][17] ), .Z(\mreg/_04366_ ) );
BUF_X1 \mreg/_12352_ ( .A(\mreg/rf[21][17] ), .Z(\mreg/_04334_ ) );
BUF_X1 \mreg/_12353_ ( .A(\mreg/rf[20][17] ), .Z(\mreg/_04302_ ) );
BUF_X1 \mreg/_12354_ ( .A(\mreg/rf[19][17] ), .Z(\mreg/_04238_ ) );
BUF_X1 \mreg/_12355_ ( .A(\mreg/rf[18][17] ), .Z(\mreg/_04206_ ) );
BUF_X1 \mreg/_12356_ ( .A(\mreg/rf[17][17] ), .Z(\mreg/_04174_ ) );
BUF_X1 \mreg/_12357_ ( .A(\mreg/rf[16][17] ), .Z(\mreg/_04142_ ) );
BUF_X1 \mreg/_12358_ ( .A(\mreg/rf[15][17] ), .Z(\mreg/_04110_ ) );
BUF_X1 \mreg/_12359_ ( .A(\mreg/rf[14][17] ), .Z(\mreg/_04078_ ) );
BUF_X1 \mreg/_12360_ ( .A(\mreg/rf[13][17] ), .Z(\mreg/_04046_ ) );
BUF_X1 \mreg/_12361_ ( .A(\mreg/rf[12][17] ), .Z(\mreg/_04014_ ) );
BUF_X1 \mreg/_12362_ ( .A(\mreg/rf[11][17] ), .Z(\mreg/_03982_ ) );
BUF_X1 \mreg/_12363_ ( .A(\mreg/rf[10][17] ), .Z(\mreg/_03950_ ) );
BUF_X1 \mreg/_12364_ ( .A(\mreg/rf[9][17] ), .Z(\mreg/_04910_ ) );
BUF_X1 \mreg/_12365_ ( .A(\mreg/rf[8][17] ), .Z(\mreg/_04878_ ) );
BUF_X1 \mreg/_12366_ ( .A(\mreg/rf[7][17] ), .Z(\mreg/_04846_ ) );
BUF_X1 \mreg/_12367_ ( .A(\mreg/rf[6][17] ), .Z(\mreg/_04814_ ) );
BUF_X1 \mreg/_12368_ ( .A(\mreg/rf[5][17] ), .Z(\mreg/_04782_ ) );
BUF_X1 \mreg/_12369_ ( .A(\mreg/rf[4][17] ), .Z(\mreg/_04750_ ) );
BUF_X1 \mreg/_12370_ ( .A(\mreg/rf[3][17] ), .Z(\mreg/_04718_ ) );
BUF_X1 \mreg/_12371_ ( .A(\mreg/rf[2][17] ), .Z(\mreg/_04622_ ) );
BUF_X1 \mreg/_12372_ ( .A(\mreg/rf[1][17] ), .Z(\mreg/_04270_ ) );
BUF_X1 \mreg/_12373_ ( .A(\mreg/_03918_ ), .Z(\mem_wdata[17] ) );
BUF_X1 \mreg/_12374_ ( .A(\mreg/_00017_ ), .Z(\mreg/_00048_ ) );
BUF_X1 \mreg/_12375_ ( .A(\mreg/rf[30][18] ), .Z(\mreg/_04655_ ) );
BUF_X1 \mreg/_12376_ ( .A(\mreg/rf[29][18] ), .Z(\mreg/_04591_ ) );
BUF_X1 \mreg/_12377_ ( .A(\mreg/rf[28][18] ), .Z(\mreg/_04559_ ) );
BUF_X1 \mreg/_12378_ ( .A(\mreg/rf[27][18] ), .Z(\mreg/_04527_ ) );
BUF_X1 \mreg/_12379_ ( .A(\mreg/rf[26][18] ), .Z(\mreg/_04495_ ) );
BUF_X1 \mreg/_12380_ ( .A(\mreg/rf[25][18] ), .Z(\mreg/_04463_ ) );
BUF_X1 \mreg/_12381_ ( .A(\mreg/rf[24][18] ), .Z(\mreg/_04431_ ) );
BUF_X1 \mreg/_12382_ ( .A(\mreg/rf[23][18] ), .Z(\mreg/_04399_ ) );
BUF_X1 \mreg/_12383_ ( .A(\mreg/rf[22][18] ), .Z(\mreg/_04367_ ) );
BUF_X1 \mreg/_12384_ ( .A(\mreg/rf[21][18] ), .Z(\mreg/_04335_ ) );
BUF_X1 \mreg/_12385_ ( .A(\mreg/rf[20][18] ), .Z(\mreg/_04303_ ) );
BUF_X1 \mreg/_12386_ ( .A(\mreg/rf[19][18] ), .Z(\mreg/_04239_ ) );
BUF_X1 \mreg/_12387_ ( .A(\mreg/rf[18][18] ), .Z(\mreg/_04207_ ) );
BUF_X1 \mreg/_12388_ ( .A(\mreg/rf[17][18] ), .Z(\mreg/_04175_ ) );
BUF_X1 \mreg/_12389_ ( .A(\mreg/rf[16][18] ), .Z(\mreg/_04143_ ) );
BUF_X1 \mreg/_12390_ ( .A(\mreg/rf[15][18] ), .Z(\mreg/_04111_ ) );
BUF_X1 \mreg/_12391_ ( .A(\mreg/rf[14][18] ), .Z(\mreg/_04079_ ) );
BUF_X1 \mreg/_12392_ ( .A(\mreg/rf[13][18] ), .Z(\mreg/_04047_ ) );
BUF_X1 \mreg/_12393_ ( .A(\mreg/rf[12][18] ), .Z(\mreg/_04015_ ) );
BUF_X1 \mreg/_12394_ ( .A(\mreg/rf[11][18] ), .Z(\mreg/_03983_ ) );
BUF_X1 \mreg/_12395_ ( .A(\mreg/rf[10][18] ), .Z(\mreg/_03951_ ) );
BUF_X1 \mreg/_12396_ ( .A(\mreg/rf[9][18] ), .Z(\mreg/_04911_ ) );
BUF_X1 \mreg/_12397_ ( .A(\mreg/rf[8][18] ), .Z(\mreg/_04879_ ) );
BUF_X1 \mreg/_12398_ ( .A(\mreg/rf[7][18] ), .Z(\mreg/_04847_ ) );
BUF_X1 \mreg/_12399_ ( .A(\mreg/rf[6][18] ), .Z(\mreg/_04815_ ) );
BUF_X1 \mreg/_12400_ ( .A(\mreg/rf[5][18] ), .Z(\mreg/_04783_ ) );
BUF_X1 \mreg/_12401_ ( .A(\mreg/rf[4][18] ), .Z(\mreg/_04751_ ) );
BUF_X1 \mreg/_12402_ ( .A(\mreg/rf[3][18] ), .Z(\mreg/_04719_ ) );
BUF_X1 \mreg/_12403_ ( .A(\mreg/rf[2][18] ), .Z(\mreg/_04623_ ) );
BUF_X1 \mreg/_12404_ ( .A(\mreg/rf[1][18] ), .Z(\mreg/_04271_ ) );
BUF_X1 \mreg/_12405_ ( .A(\mreg/_03919_ ), .Z(\mem_wdata[18] ) );
BUF_X1 \mreg/_12406_ ( .A(\mreg/_00018_ ), .Z(\mreg/_00049_ ) );
BUF_X1 \mreg/_12407_ ( .A(\mreg/rf[30][19] ), .Z(\mreg/_04656_ ) );
BUF_X1 \mreg/_12408_ ( .A(\mreg/rf[29][19] ), .Z(\mreg/_04592_ ) );
BUF_X1 \mreg/_12409_ ( .A(\mreg/rf[28][19] ), .Z(\mreg/_04560_ ) );
BUF_X1 \mreg/_12410_ ( .A(\mreg/rf[27][19] ), .Z(\mreg/_04528_ ) );
BUF_X1 \mreg/_12411_ ( .A(\mreg/rf[26][19] ), .Z(\mreg/_04496_ ) );
BUF_X1 \mreg/_12412_ ( .A(\mreg/rf[25][19] ), .Z(\mreg/_04464_ ) );
BUF_X1 \mreg/_12413_ ( .A(\mreg/rf[24][19] ), .Z(\mreg/_04432_ ) );
BUF_X1 \mreg/_12414_ ( .A(\mreg/rf[23][19] ), .Z(\mreg/_04400_ ) );
BUF_X1 \mreg/_12415_ ( .A(\mreg/rf[22][19] ), .Z(\mreg/_04368_ ) );
BUF_X1 \mreg/_12416_ ( .A(\mreg/rf[21][19] ), .Z(\mreg/_04336_ ) );
BUF_X1 \mreg/_12417_ ( .A(\mreg/rf[20][19] ), .Z(\mreg/_04304_ ) );
BUF_X1 \mreg/_12418_ ( .A(\mreg/rf[19][19] ), .Z(\mreg/_04240_ ) );
BUF_X1 \mreg/_12419_ ( .A(\mreg/rf[18][19] ), .Z(\mreg/_04208_ ) );
BUF_X1 \mreg/_12420_ ( .A(\mreg/rf[17][19] ), .Z(\mreg/_04176_ ) );
BUF_X1 \mreg/_12421_ ( .A(\mreg/rf[16][19] ), .Z(\mreg/_04144_ ) );
BUF_X1 \mreg/_12422_ ( .A(\mreg/rf[15][19] ), .Z(\mreg/_04112_ ) );
BUF_X1 \mreg/_12423_ ( .A(\mreg/rf[14][19] ), .Z(\mreg/_04080_ ) );
BUF_X1 \mreg/_12424_ ( .A(\mreg/rf[13][19] ), .Z(\mreg/_04048_ ) );
BUF_X1 \mreg/_12425_ ( .A(\mreg/rf[12][19] ), .Z(\mreg/_04016_ ) );
BUF_X1 \mreg/_12426_ ( .A(\mreg/rf[11][19] ), .Z(\mreg/_03984_ ) );
BUF_X1 \mreg/_12427_ ( .A(\mreg/rf[10][19] ), .Z(\mreg/_03952_ ) );
BUF_X1 \mreg/_12428_ ( .A(\mreg/rf[9][19] ), .Z(\mreg/_04912_ ) );
BUF_X1 \mreg/_12429_ ( .A(\mreg/rf[8][19] ), .Z(\mreg/_04880_ ) );
BUF_X1 \mreg/_12430_ ( .A(\mreg/rf[7][19] ), .Z(\mreg/_04848_ ) );
BUF_X1 \mreg/_12431_ ( .A(\mreg/rf[6][19] ), .Z(\mreg/_04816_ ) );
BUF_X1 \mreg/_12432_ ( .A(\mreg/rf[5][19] ), .Z(\mreg/_04784_ ) );
BUF_X1 \mreg/_12433_ ( .A(\mreg/rf[4][19] ), .Z(\mreg/_04752_ ) );
BUF_X1 \mreg/_12434_ ( .A(\mreg/rf[3][19] ), .Z(\mreg/_04720_ ) );
BUF_X1 \mreg/_12435_ ( .A(\mreg/rf[2][19] ), .Z(\mreg/_04624_ ) );
BUF_X1 \mreg/_12436_ ( .A(\mreg/rf[1][19] ), .Z(\mreg/_04272_ ) );
BUF_X1 \mreg/_12437_ ( .A(\mreg/_03920_ ), .Z(\mem_wdata[19] ) );
BUF_X1 \mreg/_12438_ ( .A(\mreg/_00019_ ), .Z(\mreg/_00050_ ) );
BUF_X1 \mreg/_12439_ ( .A(\mreg/rf[30][20] ), .Z(\mreg/_04658_ ) );
BUF_X1 \mreg/_12440_ ( .A(\mreg/rf[29][20] ), .Z(\mreg/_04594_ ) );
BUF_X1 \mreg/_12441_ ( .A(\mreg/rf[28][20] ), .Z(\mreg/_04562_ ) );
BUF_X1 \mreg/_12442_ ( .A(\mreg/rf[27][20] ), .Z(\mreg/_04530_ ) );
BUF_X1 \mreg/_12443_ ( .A(\mreg/rf[26][20] ), .Z(\mreg/_04498_ ) );
BUF_X1 \mreg/_12444_ ( .A(\mreg/rf[25][20] ), .Z(\mreg/_04466_ ) );
BUF_X1 \mreg/_12445_ ( .A(\mreg/rf[24][20] ), .Z(\mreg/_04434_ ) );
BUF_X1 \mreg/_12446_ ( .A(\mreg/rf[23][20] ), .Z(\mreg/_04402_ ) );
BUF_X1 \mreg/_12447_ ( .A(\mreg/rf[22][20] ), .Z(\mreg/_04370_ ) );
BUF_X1 \mreg/_12448_ ( .A(\mreg/rf[21][20] ), .Z(\mreg/_04338_ ) );
BUF_X1 \mreg/_12449_ ( .A(\mreg/rf[20][20] ), .Z(\mreg/_04306_ ) );
BUF_X1 \mreg/_12450_ ( .A(\mreg/rf[19][20] ), .Z(\mreg/_04242_ ) );
BUF_X1 \mreg/_12451_ ( .A(\mreg/rf[18][20] ), .Z(\mreg/_04210_ ) );
BUF_X1 \mreg/_12452_ ( .A(\mreg/rf[17][20] ), .Z(\mreg/_04178_ ) );
BUF_X1 \mreg/_12453_ ( .A(\mreg/rf[16][20] ), .Z(\mreg/_04146_ ) );
BUF_X1 \mreg/_12454_ ( .A(\mreg/rf[15][20] ), .Z(\mreg/_04114_ ) );
BUF_X1 \mreg/_12455_ ( .A(\mreg/rf[14][20] ), .Z(\mreg/_04082_ ) );
BUF_X1 \mreg/_12456_ ( .A(\mreg/rf[13][20] ), .Z(\mreg/_04050_ ) );
BUF_X1 \mreg/_12457_ ( .A(\mreg/rf[12][20] ), .Z(\mreg/_04018_ ) );
BUF_X1 \mreg/_12458_ ( .A(\mreg/rf[11][20] ), .Z(\mreg/_03986_ ) );
BUF_X1 \mreg/_12459_ ( .A(\mreg/rf[10][20] ), .Z(\mreg/_03954_ ) );
BUF_X1 \mreg/_12460_ ( .A(\mreg/rf[9][20] ), .Z(\mreg/_04914_ ) );
BUF_X1 \mreg/_12461_ ( .A(\mreg/rf[8][20] ), .Z(\mreg/_04882_ ) );
BUF_X1 \mreg/_12462_ ( .A(\mreg/rf[7][20] ), .Z(\mreg/_04850_ ) );
BUF_X1 \mreg/_12463_ ( .A(\mreg/rf[6][20] ), .Z(\mreg/_04818_ ) );
BUF_X1 \mreg/_12464_ ( .A(\mreg/rf[5][20] ), .Z(\mreg/_04786_ ) );
BUF_X1 \mreg/_12465_ ( .A(\mreg/rf[4][20] ), .Z(\mreg/_04754_ ) );
BUF_X1 \mreg/_12466_ ( .A(\mreg/rf[3][20] ), .Z(\mreg/_04722_ ) );
BUF_X1 \mreg/_12467_ ( .A(\mreg/rf[2][20] ), .Z(\mreg/_04626_ ) );
BUF_X1 \mreg/_12468_ ( .A(\mreg/rf[1][20] ), .Z(\mreg/_04274_ ) );
BUF_X1 \mreg/_12469_ ( .A(\mreg/_03922_ ), .Z(\mem_wdata[20] ) );
BUF_X1 \mreg/_12470_ ( .A(\mreg/_00020_ ), .Z(\mreg/_00051_ ) );
BUF_X1 \mreg/_12471_ ( .A(\mreg/rf[30][21] ), .Z(\mreg/_04659_ ) );
BUF_X1 \mreg/_12472_ ( .A(\mreg/rf[29][21] ), .Z(\mreg/_04595_ ) );
BUF_X1 \mreg/_12473_ ( .A(\mreg/rf[28][21] ), .Z(\mreg/_04563_ ) );
BUF_X1 \mreg/_12474_ ( .A(\mreg/rf[27][21] ), .Z(\mreg/_04531_ ) );
BUF_X1 \mreg/_12475_ ( .A(\mreg/rf[26][21] ), .Z(\mreg/_04499_ ) );
BUF_X1 \mreg/_12476_ ( .A(\mreg/rf[25][21] ), .Z(\mreg/_04467_ ) );
BUF_X1 \mreg/_12477_ ( .A(\mreg/rf[24][21] ), .Z(\mreg/_04435_ ) );
BUF_X1 \mreg/_12478_ ( .A(\mreg/rf[23][21] ), .Z(\mreg/_04403_ ) );
BUF_X1 \mreg/_12479_ ( .A(\mreg/rf[22][21] ), .Z(\mreg/_04371_ ) );
BUF_X1 \mreg/_12480_ ( .A(\mreg/rf[21][21] ), .Z(\mreg/_04339_ ) );
BUF_X1 \mreg/_12481_ ( .A(\mreg/rf[20][21] ), .Z(\mreg/_04307_ ) );
BUF_X1 \mreg/_12482_ ( .A(\mreg/rf[19][21] ), .Z(\mreg/_04243_ ) );
BUF_X1 \mreg/_12483_ ( .A(\mreg/rf[18][21] ), .Z(\mreg/_04211_ ) );
BUF_X1 \mreg/_12484_ ( .A(\mreg/rf[17][21] ), .Z(\mreg/_04179_ ) );
BUF_X1 \mreg/_12485_ ( .A(\mreg/rf[16][21] ), .Z(\mreg/_04147_ ) );
BUF_X1 \mreg/_12486_ ( .A(\mreg/rf[15][21] ), .Z(\mreg/_04115_ ) );
BUF_X1 \mreg/_12487_ ( .A(\mreg/rf[14][21] ), .Z(\mreg/_04083_ ) );
BUF_X1 \mreg/_12488_ ( .A(\mreg/rf[13][21] ), .Z(\mreg/_04051_ ) );
BUF_X1 \mreg/_12489_ ( .A(\mreg/rf[12][21] ), .Z(\mreg/_04019_ ) );
BUF_X1 \mreg/_12490_ ( .A(\mreg/rf[11][21] ), .Z(\mreg/_03987_ ) );
BUF_X1 \mreg/_12491_ ( .A(\mreg/rf[10][21] ), .Z(\mreg/_03955_ ) );
BUF_X1 \mreg/_12492_ ( .A(\mreg/rf[9][21] ), .Z(\mreg/_04915_ ) );
BUF_X1 \mreg/_12493_ ( .A(\mreg/rf[8][21] ), .Z(\mreg/_04883_ ) );
BUF_X1 \mreg/_12494_ ( .A(\mreg/rf[7][21] ), .Z(\mreg/_04851_ ) );
BUF_X1 \mreg/_12495_ ( .A(\mreg/rf[6][21] ), .Z(\mreg/_04819_ ) );
BUF_X1 \mreg/_12496_ ( .A(\mreg/rf[5][21] ), .Z(\mreg/_04787_ ) );
BUF_X1 \mreg/_12497_ ( .A(\mreg/rf[4][21] ), .Z(\mreg/_04755_ ) );
BUF_X1 \mreg/_12498_ ( .A(\mreg/rf[3][21] ), .Z(\mreg/_04723_ ) );
BUF_X1 \mreg/_12499_ ( .A(\mreg/rf[2][21] ), .Z(\mreg/_04627_ ) );
BUF_X1 \mreg/_12500_ ( .A(\mreg/rf[1][21] ), .Z(\mreg/_04275_ ) );
BUF_X1 \mreg/_12501_ ( .A(\mreg/_03923_ ), .Z(\mem_wdata[21] ) );
BUF_X1 \mreg/_12502_ ( .A(\mreg/_00021_ ), .Z(\mreg/_00052_ ) );
BUF_X1 \mreg/_12503_ ( .A(\mreg/rf[30][22] ), .Z(\mreg/_04660_ ) );
BUF_X1 \mreg/_12504_ ( .A(\mreg/rf[29][22] ), .Z(\mreg/_04596_ ) );
BUF_X1 \mreg/_12505_ ( .A(\mreg/rf[28][22] ), .Z(\mreg/_04564_ ) );
BUF_X1 \mreg/_12506_ ( .A(\mreg/rf[27][22] ), .Z(\mreg/_04532_ ) );
BUF_X1 \mreg/_12507_ ( .A(\mreg/rf[26][22] ), .Z(\mreg/_04500_ ) );
BUF_X1 \mreg/_12508_ ( .A(\mreg/rf[25][22] ), .Z(\mreg/_04468_ ) );
BUF_X1 \mreg/_12509_ ( .A(\mreg/rf[24][22] ), .Z(\mreg/_04436_ ) );
BUF_X1 \mreg/_12510_ ( .A(\mreg/rf[23][22] ), .Z(\mreg/_04404_ ) );
BUF_X1 \mreg/_12511_ ( .A(\mreg/rf[22][22] ), .Z(\mreg/_04372_ ) );
BUF_X1 \mreg/_12512_ ( .A(\mreg/rf[21][22] ), .Z(\mreg/_04340_ ) );
BUF_X1 \mreg/_12513_ ( .A(\mreg/rf[20][22] ), .Z(\mreg/_04308_ ) );
BUF_X1 \mreg/_12514_ ( .A(\mreg/rf[19][22] ), .Z(\mreg/_04244_ ) );
BUF_X1 \mreg/_12515_ ( .A(\mreg/rf[18][22] ), .Z(\mreg/_04212_ ) );
BUF_X1 \mreg/_12516_ ( .A(\mreg/rf[17][22] ), .Z(\mreg/_04180_ ) );
BUF_X1 \mreg/_12517_ ( .A(\mreg/rf[16][22] ), .Z(\mreg/_04148_ ) );
BUF_X1 \mreg/_12518_ ( .A(\mreg/rf[15][22] ), .Z(\mreg/_04116_ ) );
BUF_X1 \mreg/_12519_ ( .A(\mreg/rf[14][22] ), .Z(\mreg/_04084_ ) );
BUF_X1 \mreg/_12520_ ( .A(\mreg/rf[13][22] ), .Z(\mreg/_04052_ ) );
BUF_X1 \mreg/_12521_ ( .A(\mreg/rf[12][22] ), .Z(\mreg/_04020_ ) );
BUF_X1 \mreg/_12522_ ( .A(\mreg/rf[11][22] ), .Z(\mreg/_03988_ ) );
BUF_X1 \mreg/_12523_ ( .A(\mreg/rf[10][22] ), .Z(\mreg/_03956_ ) );
BUF_X1 \mreg/_12524_ ( .A(\mreg/rf[9][22] ), .Z(\mreg/_04916_ ) );
BUF_X1 \mreg/_12525_ ( .A(\mreg/rf[8][22] ), .Z(\mreg/_04884_ ) );
BUF_X1 \mreg/_12526_ ( .A(\mreg/rf[7][22] ), .Z(\mreg/_04852_ ) );
BUF_X1 \mreg/_12527_ ( .A(\mreg/rf[6][22] ), .Z(\mreg/_04820_ ) );
BUF_X1 \mreg/_12528_ ( .A(\mreg/rf[5][22] ), .Z(\mreg/_04788_ ) );
BUF_X1 \mreg/_12529_ ( .A(\mreg/rf[4][22] ), .Z(\mreg/_04756_ ) );
BUF_X1 \mreg/_12530_ ( .A(\mreg/rf[3][22] ), .Z(\mreg/_04724_ ) );
BUF_X1 \mreg/_12531_ ( .A(\mreg/rf[2][22] ), .Z(\mreg/_04628_ ) );
BUF_X1 \mreg/_12532_ ( .A(\mreg/rf[1][22] ), .Z(\mreg/_04276_ ) );
BUF_X1 \mreg/_12533_ ( .A(\mreg/_03924_ ), .Z(\mem_wdata[22] ) );
BUF_X1 \mreg/_12534_ ( .A(\mreg/_00022_ ), .Z(\mreg/_00053_ ) );
BUF_X1 \mreg/_12535_ ( .A(\mreg/rf[30][23] ), .Z(\mreg/_04661_ ) );
BUF_X1 \mreg/_12536_ ( .A(\mreg/rf[29][23] ), .Z(\mreg/_04597_ ) );
BUF_X1 \mreg/_12537_ ( .A(\mreg/rf[28][23] ), .Z(\mreg/_04565_ ) );
BUF_X1 \mreg/_12538_ ( .A(\mreg/rf[27][23] ), .Z(\mreg/_04533_ ) );
BUF_X1 \mreg/_12539_ ( .A(\mreg/rf[26][23] ), .Z(\mreg/_04501_ ) );
BUF_X1 \mreg/_12540_ ( .A(\mreg/rf[25][23] ), .Z(\mreg/_04469_ ) );
BUF_X1 \mreg/_12541_ ( .A(\mreg/rf[24][23] ), .Z(\mreg/_04437_ ) );
BUF_X1 \mreg/_12542_ ( .A(\mreg/rf[23][23] ), .Z(\mreg/_04405_ ) );
BUF_X1 \mreg/_12543_ ( .A(\mreg/rf[22][23] ), .Z(\mreg/_04373_ ) );
BUF_X1 \mreg/_12544_ ( .A(\mreg/rf[21][23] ), .Z(\mreg/_04341_ ) );
BUF_X1 \mreg/_12545_ ( .A(\mreg/rf[20][23] ), .Z(\mreg/_04309_ ) );
BUF_X1 \mreg/_12546_ ( .A(\mreg/rf[19][23] ), .Z(\mreg/_04245_ ) );
BUF_X1 \mreg/_12547_ ( .A(\mreg/rf[18][23] ), .Z(\mreg/_04213_ ) );
BUF_X1 \mreg/_12548_ ( .A(\mreg/rf[17][23] ), .Z(\mreg/_04181_ ) );
BUF_X1 \mreg/_12549_ ( .A(\mreg/rf[16][23] ), .Z(\mreg/_04149_ ) );
BUF_X1 \mreg/_12550_ ( .A(\mreg/rf[15][23] ), .Z(\mreg/_04117_ ) );
BUF_X1 \mreg/_12551_ ( .A(\mreg/rf[14][23] ), .Z(\mreg/_04085_ ) );
BUF_X1 \mreg/_12552_ ( .A(\mreg/rf[13][23] ), .Z(\mreg/_04053_ ) );
BUF_X1 \mreg/_12553_ ( .A(\mreg/rf[12][23] ), .Z(\mreg/_04021_ ) );
BUF_X1 \mreg/_12554_ ( .A(\mreg/rf[11][23] ), .Z(\mreg/_03989_ ) );
BUF_X1 \mreg/_12555_ ( .A(\mreg/rf[10][23] ), .Z(\mreg/_03957_ ) );
BUF_X1 \mreg/_12556_ ( .A(\mreg/rf[9][23] ), .Z(\mreg/_04917_ ) );
BUF_X1 \mreg/_12557_ ( .A(\mreg/rf[8][23] ), .Z(\mreg/_04885_ ) );
BUF_X1 \mreg/_12558_ ( .A(\mreg/rf[7][23] ), .Z(\mreg/_04853_ ) );
BUF_X1 \mreg/_12559_ ( .A(\mreg/rf[6][23] ), .Z(\mreg/_04821_ ) );
BUF_X1 \mreg/_12560_ ( .A(\mreg/rf[5][23] ), .Z(\mreg/_04789_ ) );
BUF_X1 \mreg/_12561_ ( .A(\mreg/rf[4][23] ), .Z(\mreg/_04757_ ) );
BUF_X1 \mreg/_12562_ ( .A(\mreg/rf[3][23] ), .Z(\mreg/_04725_ ) );
BUF_X1 \mreg/_12563_ ( .A(\mreg/rf[2][23] ), .Z(\mreg/_04629_ ) );
BUF_X1 \mreg/_12564_ ( .A(\mreg/rf[1][23] ), .Z(\mreg/_04277_ ) );
BUF_X1 \mreg/_12565_ ( .A(\mreg/_03925_ ), .Z(\mem_wdata[23] ) );
BUF_X1 \mreg/_12566_ ( .A(\mreg/_00023_ ), .Z(\mreg/_00054_ ) );
BUF_X1 \mreg/_12567_ ( .A(\mreg/rf[30][24] ), .Z(\mreg/_04662_ ) );
BUF_X1 \mreg/_12568_ ( .A(\mreg/rf[29][24] ), .Z(\mreg/_04598_ ) );
BUF_X1 \mreg/_12569_ ( .A(\mreg/rf[28][24] ), .Z(\mreg/_04566_ ) );
BUF_X1 \mreg/_12570_ ( .A(\mreg/rf[27][24] ), .Z(\mreg/_04534_ ) );
BUF_X1 \mreg/_12571_ ( .A(\mreg/rf[26][24] ), .Z(\mreg/_04502_ ) );
BUF_X1 \mreg/_12572_ ( .A(\mreg/rf[25][24] ), .Z(\mreg/_04470_ ) );
BUF_X1 \mreg/_12573_ ( .A(\mreg/rf[24][24] ), .Z(\mreg/_04438_ ) );
BUF_X1 \mreg/_12574_ ( .A(\mreg/rf[23][24] ), .Z(\mreg/_04406_ ) );
BUF_X1 \mreg/_12575_ ( .A(\mreg/rf[22][24] ), .Z(\mreg/_04374_ ) );
BUF_X1 \mreg/_12576_ ( .A(\mreg/rf[21][24] ), .Z(\mreg/_04342_ ) );
BUF_X1 \mreg/_12577_ ( .A(\mreg/rf[20][24] ), .Z(\mreg/_04310_ ) );
BUF_X1 \mreg/_12578_ ( .A(\mreg/rf[19][24] ), .Z(\mreg/_04246_ ) );
BUF_X1 \mreg/_12579_ ( .A(\mreg/rf[18][24] ), .Z(\mreg/_04214_ ) );
BUF_X1 \mreg/_12580_ ( .A(\mreg/rf[17][24] ), .Z(\mreg/_04182_ ) );
BUF_X1 \mreg/_12581_ ( .A(\mreg/rf[16][24] ), .Z(\mreg/_04150_ ) );
BUF_X1 \mreg/_12582_ ( .A(\mreg/rf[15][24] ), .Z(\mreg/_04118_ ) );
BUF_X1 \mreg/_12583_ ( .A(\mreg/rf[14][24] ), .Z(\mreg/_04086_ ) );
BUF_X1 \mreg/_12584_ ( .A(\mreg/rf[13][24] ), .Z(\mreg/_04054_ ) );
BUF_X1 \mreg/_12585_ ( .A(\mreg/rf[12][24] ), .Z(\mreg/_04022_ ) );
BUF_X1 \mreg/_12586_ ( .A(\mreg/rf[11][24] ), .Z(\mreg/_03990_ ) );
BUF_X1 \mreg/_12587_ ( .A(\mreg/rf[10][24] ), .Z(\mreg/_03958_ ) );
BUF_X1 \mreg/_12588_ ( .A(\mreg/rf[9][24] ), .Z(\mreg/_04918_ ) );
BUF_X1 \mreg/_12589_ ( .A(\mreg/rf[8][24] ), .Z(\mreg/_04886_ ) );
BUF_X1 \mreg/_12590_ ( .A(\mreg/rf[7][24] ), .Z(\mreg/_04854_ ) );
BUF_X1 \mreg/_12591_ ( .A(\mreg/rf[6][24] ), .Z(\mreg/_04822_ ) );
BUF_X1 \mreg/_12592_ ( .A(\mreg/rf[5][24] ), .Z(\mreg/_04790_ ) );
BUF_X1 \mreg/_12593_ ( .A(\mreg/rf[4][24] ), .Z(\mreg/_04758_ ) );
BUF_X1 \mreg/_12594_ ( .A(\mreg/rf[3][24] ), .Z(\mreg/_04726_ ) );
BUF_X1 \mreg/_12595_ ( .A(\mreg/rf[2][24] ), .Z(\mreg/_04630_ ) );
BUF_X1 \mreg/_12596_ ( .A(\mreg/rf[1][24] ), .Z(\mreg/_04278_ ) );
BUF_X1 \mreg/_12597_ ( .A(\mreg/_03926_ ), .Z(\mem_wdata[24] ) );
BUF_X1 \mreg/_12598_ ( .A(\mreg/_00024_ ), .Z(\mreg/_00055_ ) );
BUF_X1 \mreg/_12599_ ( .A(\mreg/rf[30][25] ), .Z(\mreg/_04663_ ) );
BUF_X1 \mreg/_12600_ ( .A(\mreg/rf[29][25] ), .Z(\mreg/_04599_ ) );
BUF_X1 \mreg/_12601_ ( .A(\mreg/rf[28][25] ), .Z(\mreg/_04567_ ) );
BUF_X1 \mreg/_12602_ ( .A(\mreg/rf[27][25] ), .Z(\mreg/_04535_ ) );
BUF_X1 \mreg/_12603_ ( .A(\mreg/rf[26][25] ), .Z(\mreg/_04503_ ) );
BUF_X1 \mreg/_12604_ ( .A(\mreg/rf[25][25] ), .Z(\mreg/_04471_ ) );
BUF_X1 \mreg/_12605_ ( .A(\mreg/rf[24][25] ), .Z(\mreg/_04439_ ) );
BUF_X1 \mreg/_12606_ ( .A(\mreg/rf[23][25] ), .Z(\mreg/_04407_ ) );
BUF_X1 \mreg/_12607_ ( .A(\mreg/rf[22][25] ), .Z(\mreg/_04375_ ) );
BUF_X1 \mreg/_12608_ ( .A(\mreg/rf[21][25] ), .Z(\mreg/_04343_ ) );
BUF_X1 \mreg/_12609_ ( .A(\mreg/rf[20][25] ), .Z(\mreg/_04311_ ) );
BUF_X1 \mreg/_12610_ ( .A(\mreg/rf[19][25] ), .Z(\mreg/_04247_ ) );
BUF_X1 \mreg/_12611_ ( .A(\mreg/rf[18][25] ), .Z(\mreg/_04215_ ) );
BUF_X1 \mreg/_12612_ ( .A(\mreg/rf[17][25] ), .Z(\mreg/_04183_ ) );
BUF_X1 \mreg/_12613_ ( .A(\mreg/rf[16][25] ), .Z(\mreg/_04151_ ) );
BUF_X1 \mreg/_12614_ ( .A(\mreg/rf[15][25] ), .Z(\mreg/_04119_ ) );
BUF_X1 \mreg/_12615_ ( .A(\mreg/rf[14][25] ), .Z(\mreg/_04087_ ) );
BUF_X1 \mreg/_12616_ ( .A(\mreg/rf[13][25] ), .Z(\mreg/_04055_ ) );
BUF_X1 \mreg/_12617_ ( .A(\mreg/rf[12][25] ), .Z(\mreg/_04023_ ) );
BUF_X1 \mreg/_12618_ ( .A(\mreg/rf[11][25] ), .Z(\mreg/_03991_ ) );
BUF_X1 \mreg/_12619_ ( .A(\mreg/rf[10][25] ), .Z(\mreg/_03959_ ) );
BUF_X1 \mreg/_12620_ ( .A(\mreg/rf[9][25] ), .Z(\mreg/_04919_ ) );
BUF_X1 \mreg/_12621_ ( .A(\mreg/rf[8][25] ), .Z(\mreg/_04887_ ) );
BUF_X1 \mreg/_12622_ ( .A(\mreg/rf[7][25] ), .Z(\mreg/_04855_ ) );
BUF_X1 \mreg/_12623_ ( .A(\mreg/rf[6][25] ), .Z(\mreg/_04823_ ) );
BUF_X1 \mreg/_12624_ ( .A(\mreg/rf[5][25] ), .Z(\mreg/_04791_ ) );
BUF_X1 \mreg/_12625_ ( .A(\mreg/rf[4][25] ), .Z(\mreg/_04759_ ) );
BUF_X1 \mreg/_12626_ ( .A(\mreg/rf[3][25] ), .Z(\mreg/_04727_ ) );
BUF_X1 \mreg/_12627_ ( .A(\mreg/rf[2][25] ), .Z(\mreg/_04631_ ) );
BUF_X1 \mreg/_12628_ ( .A(\mreg/rf[1][25] ), .Z(\mreg/_04279_ ) );
BUF_X1 \mreg/_12629_ ( .A(\mreg/_03927_ ), .Z(\mem_wdata[25] ) );
BUF_X1 \mreg/_12630_ ( .A(\mreg/_00025_ ), .Z(\mreg/_00056_ ) );
BUF_X1 \mreg/_12631_ ( .A(\mreg/rf[30][26] ), .Z(\mreg/_04664_ ) );
BUF_X1 \mreg/_12632_ ( .A(\mreg/rf[29][26] ), .Z(\mreg/_04600_ ) );
BUF_X1 \mreg/_12633_ ( .A(\mreg/rf[28][26] ), .Z(\mreg/_04568_ ) );
BUF_X1 \mreg/_12634_ ( .A(\mreg/rf[27][26] ), .Z(\mreg/_04536_ ) );
BUF_X1 \mreg/_12635_ ( .A(\mreg/rf[26][26] ), .Z(\mreg/_04504_ ) );
BUF_X1 \mreg/_12636_ ( .A(\mreg/rf[25][26] ), .Z(\mreg/_04472_ ) );
BUF_X1 \mreg/_12637_ ( .A(\mreg/rf[24][26] ), .Z(\mreg/_04440_ ) );
BUF_X1 \mreg/_12638_ ( .A(\mreg/rf[23][26] ), .Z(\mreg/_04408_ ) );
BUF_X1 \mreg/_12639_ ( .A(\mreg/rf[22][26] ), .Z(\mreg/_04376_ ) );
BUF_X1 \mreg/_12640_ ( .A(\mreg/rf[21][26] ), .Z(\mreg/_04344_ ) );
BUF_X1 \mreg/_12641_ ( .A(\mreg/rf[20][26] ), .Z(\mreg/_04312_ ) );
BUF_X1 \mreg/_12642_ ( .A(\mreg/rf[19][26] ), .Z(\mreg/_04248_ ) );
BUF_X1 \mreg/_12643_ ( .A(\mreg/rf[18][26] ), .Z(\mreg/_04216_ ) );
BUF_X1 \mreg/_12644_ ( .A(\mreg/rf[17][26] ), .Z(\mreg/_04184_ ) );
BUF_X1 \mreg/_12645_ ( .A(\mreg/rf[16][26] ), .Z(\mreg/_04152_ ) );
BUF_X1 \mreg/_12646_ ( .A(\mreg/rf[15][26] ), .Z(\mreg/_04120_ ) );
BUF_X1 \mreg/_12647_ ( .A(\mreg/rf[14][26] ), .Z(\mreg/_04088_ ) );
BUF_X1 \mreg/_12648_ ( .A(\mreg/rf[13][26] ), .Z(\mreg/_04056_ ) );
BUF_X1 \mreg/_12649_ ( .A(\mreg/rf[12][26] ), .Z(\mreg/_04024_ ) );
BUF_X1 \mreg/_12650_ ( .A(\mreg/rf[11][26] ), .Z(\mreg/_03992_ ) );
BUF_X1 \mreg/_12651_ ( .A(\mreg/rf[10][26] ), .Z(\mreg/_03960_ ) );
BUF_X1 \mreg/_12652_ ( .A(\mreg/rf[9][26] ), .Z(\mreg/_04920_ ) );
BUF_X1 \mreg/_12653_ ( .A(\mreg/rf[8][26] ), .Z(\mreg/_04888_ ) );
BUF_X1 \mreg/_12654_ ( .A(\mreg/rf[7][26] ), .Z(\mreg/_04856_ ) );
BUF_X1 \mreg/_12655_ ( .A(\mreg/rf[6][26] ), .Z(\mreg/_04824_ ) );
BUF_X1 \mreg/_12656_ ( .A(\mreg/rf[5][26] ), .Z(\mreg/_04792_ ) );
BUF_X1 \mreg/_12657_ ( .A(\mreg/rf[4][26] ), .Z(\mreg/_04760_ ) );
BUF_X1 \mreg/_12658_ ( .A(\mreg/rf[3][26] ), .Z(\mreg/_04728_ ) );
BUF_X1 \mreg/_12659_ ( .A(\mreg/rf[2][26] ), .Z(\mreg/_04632_ ) );
BUF_X1 \mreg/_12660_ ( .A(\mreg/rf[1][26] ), .Z(\mreg/_04280_ ) );
BUF_X1 \mreg/_12661_ ( .A(\mreg/_03928_ ), .Z(\mem_wdata[26] ) );
BUF_X1 \mreg/_12662_ ( .A(\mreg/_00026_ ), .Z(\mreg/_00057_ ) );
BUF_X1 \mreg/_12663_ ( .A(\mreg/rf[30][27] ), .Z(\mreg/_04665_ ) );
BUF_X1 \mreg/_12664_ ( .A(\mreg/rf[29][27] ), .Z(\mreg/_04601_ ) );
BUF_X1 \mreg/_12665_ ( .A(\mreg/rf[28][27] ), .Z(\mreg/_04569_ ) );
BUF_X1 \mreg/_12666_ ( .A(\mreg/rf[27][27] ), .Z(\mreg/_04537_ ) );
BUF_X1 \mreg/_12667_ ( .A(\mreg/rf[26][27] ), .Z(\mreg/_04505_ ) );
BUF_X1 \mreg/_12668_ ( .A(\mreg/rf[25][27] ), .Z(\mreg/_04473_ ) );
BUF_X1 \mreg/_12669_ ( .A(\mreg/rf[24][27] ), .Z(\mreg/_04441_ ) );
BUF_X1 \mreg/_12670_ ( .A(\mreg/rf[23][27] ), .Z(\mreg/_04409_ ) );
BUF_X1 \mreg/_12671_ ( .A(\mreg/rf[22][27] ), .Z(\mreg/_04377_ ) );
BUF_X1 \mreg/_12672_ ( .A(\mreg/rf[21][27] ), .Z(\mreg/_04345_ ) );
BUF_X1 \mreg/_12673_ ( .A(\mreg/rf[20][27] ), .Z(\mreg/_04313_ ) );
BUF_X1 \mreg/_12674_ ( .A(\mreg/rf[19][27] ), .Z(\mreg/_04249_ ) );
BUF_X1 \mreg/_12675_ ( .A(\mreg/rf[18][27] ), .Z(\mreg/_04217_ ) );
BUF_X1 \mreg/_12676_ ( .A(\mreg/rf[17][27] ), .Z(\mreg/_04185_ ) );
BUF_X1 \mreg/_12677_ ( .A(\mreg/rf[16][27] ), .Z(\mreg/_04153_ ) );
BUF_X1 \mreg/_12678_ ( .A(\mreg/rf[15][27] ), .Z(\mreg/_04121_ ) );
BUF_X1 \mreg/_12679_ ( .A(\mreg/rf[14][27] ), .Z(\mreg/_04089_ ) );
BUF_X1 \mreg/_12680_ ( .A(\mreg/rf[13][27] ), .Z(\mreg/_04057_ ) );
BUF_X1 \mreg/_12681_ ( .A(\mreg/rf[12][27] ), .Z(\mreg/_04025_ ) );
BUF_X1 \mreg/_12682_ ( .A(\mreg/rf[11][27] ), .Z(\mreg/_03993_ ) );
BUF_X1 \mreg/_12683_ ( .A(\mreg/rf[10][27] ), .Z(\mreg/_03961_ ) );
BUF_X1 \mreg/_12684_ ( .A(\mreg/rf[9][27] ), .Z(\mreg/_04921_ ) );
BUF_X1 \mreg/_12685_ ( .A(\mreg/rf[8][27] ), .Z(\mreg/_04889_ ) );
BUF_X1 \mreg/_12686_ ( .A(\mreg/rf[7][27] ), .Z(\mreg/_04857_ ) );
BUF_X1 \mreg/_12687_ ( .A(\mreg/rf[6][27] ), .Z(\mreg/_04825_ ) );
BUF_X1 \mreg/_12688_ ( .A(\mreg/rf[5][27] ), .Z(\mreg/_04793_ ) );
BUF_X1 \mreg/_12689_ ( .A(\mreg/rf[4][27] ), .Z(\mreg/_04761_ ) );
BUF_X1 \mreg/_12690_ ( .A(\mreg/rf[3][27] ), .Z(\mreg/_04729_ ) );
BUF_X1 \mreg/_12691_ ( .A(\mreg/rf[2][27] ), .Z(\mreg/_04633_ ) );
BUF_X1 \mreg/_12692_ ( .A(\mreg/rf[1][27] ), .Z(\mreg/_04281_ ) );
BUF_X1 \mreg/_12693_ ( .A(\mreg/_03929_ ), .Z(\mem_wdata[27] ) );
BUF_X1 \mreg/_12694_ ( .A(\mreg/_00027_ ), .Z(\mreg/_00058_ ) );
BUF_X1 \mreg/_12695_ ( .A(\mreg/rf[30][28] ), .Z(\mreg/_04666_ ) );
BUF_X1 \mreg/_12696_ ( .A(\mreg/rf[29][28] ), .Z(\mreg/_04602_ ) );
BUF_X1 \mreg/_12697_ ( .A(\mreg/rf[28][28] ), .Z(\mreg/_04570_ ) );
BUF_X1 \mreg/_12698_ ( .A(\mreg/rf[27][28] ), .Z(\mreg/_04538_ ) );
BUF_X1 \mreg/_12699_ ( .A(\mreg/rf[26][28] ), .Z(\mreg/_04506_ ) );
BUF_X1 \mreg/_12700_ ( .A(\mreg/rf[25][28] ), .Z(\mreg/_04474_ ) );
BUF_X1 \mreg/_12701_ ( .A(\mreg/rf[24][28] ), .Z(\mreg/_04442_ ) );
BUF_X1 \mreg/_12702_ ( .A(\mreg/rf[23][28] ), .Z(\mreg/_04410_ ) );
BUF_X1 \mreg/_12703_ ( .A(\mreg/rf[22][28] ), .Z(\mreg/_04378_ ) );
BUF_X1 \mreg/_12704_ ( .A(\mreg/rf[21][28] ), .Z(\mreg/_04346_ ) );
BUF_X1 \mreg/_12705_ ( .A(\mreg/rf[20][28] ), .Z(\mreg/_04314_ ) );
BUF_X1 \mreg/_12706_ ( .A(\mreg/rf[19][28] ), .Z(\mreg/_04250_ ) );
BUF_X1 \mreg/_12707_ ( .A(\mreg/rf[18][28] ), .Z(\mreg/_04218_ ) );
BUF_X1 \mreg/_12708_ ( .A(\mreg/rf[17][28] ), .Z(\mreg/_04186_ ) );
BUF_X1 \mreg/_12709_ ( .A(\mreg/rf[16][28] ), .Z(\mreg/_04154_ ) );
BUF_X1 \mreg/_12710_ ( .A(\mreg/rf[15][28] ), .Z(\mreg/_04122_ ) );
BUF_X1 \mreg/_12711_ ( .A(\mreg/rf[14][28] ), .Z(\mreg/_04090_ ) );
BUF_X1 \mreg/_12712_ ( .A(\mreg/rf[13][28] ), .Z(\mreg/_04058_ ) );
BUF_X1 \mreg/_12713_ ( .A(\mreg/rf[12][28] ), .Z(\mreg/_04026_ ) );
BUF_X1 \mreg/_12714_ ( .A(\mreg/rf[11][28] ), .Z(\mreg/_03994_ ) );
BUF_X1 \mreg/_12715_ ( .A(\mreg/rf[10][28] ), .Z(\mreg/_03962_ ) );
BUF_X1 \mreg/_12716_ ( .A(\mreg/rf[9][28] ), .Z(\mreg/_04922_ ) );
BUF_X1 \mreg/_12717_ ( .A(\mreg/rf[8][28] ), .Z(\mreg/_04890_ ) );
BUF_X1 \mreg/_12718_ ( .A(\mreg/rf[7][28] ), .Z(\mreg/_04858_ ) );
BUF_X1 \mreg/_12719_ ( .A(\mreg/rf[6][28] ), .Z(\mreg/_04826_ ) );
BUF_X1 \mreg/_12720_ ( .A(\mreg/rf[5][28] ), .Z(\mreg/_04794_ ) );
BUF_X1 \mreg/_12721_ ( .A(\mreg/rf[4][28] ), .Z(\mreg/_04762_ ) );
BUF_X1 \mreg/_12722_ ( .A(\mreg/rf[3][28] ), .Z(\mreg/_04730_ ) );
BUF_X1 \mreg/_12723_ ( .A(\mreg/rf[2][28] ), .Z(\mreg/_04634_ ) );
BUF_X1 \mreg/_12724_ ( .A(\mreg/rf[1][28] ), .Z(\mreg/_04282_ ) );
BUF_X1 \mreg/_12725_ ( .A(\mreg/_03930_ ), .Z(\mem_wdata[28] ) );
BUF_X1 \mreg/_12726_ ( .A(\mreg/_00028_ ), .Z(\mreg/_00059_ ) );
BUF_X1 \mreg/_12727_ ( .A(\mreg/rf[30][29] ), .Z(\mreg/_04667_ ) );
BUF_X1 \mreg/_12728_ ( .A(\mreg/rf[29][29] ), .Z(\mreg/_04603_ ) );
BUF_X1 \mreg/_12729_ ( .A(\mreg/rf[28][29] ), .Z(\mreg/_04571_ ) );
BUF_X1 \mreg/_12730_ ( .A(\mreg/rf[27][29] ), .Z(\mreg/_04539_ ) );
BUF_X1 \mreg/_12731_ ( .A(\mreg/rf[26][29] ), .Z(\mreg/_04507_ ) );
BUF_X1 \mreg/_12732_ ( .A(\mreg/rf[25][29] ), .Z(\mreg/_04475_ ) );
BUF_X1 \mreg/_12733_ ( .A(\mreg/rf[24][29] ), .Z(\mreg/_04443_ ) );
BUF_X1 \mreg/_12734_ ( .A(\mreg/rf[23][29] ), .Z(\mreg/_04411_ ) );
BUF_X1 \mreg/_12735_ ( .A(\mreg/rf[22][29] ), .Z(\mreg/_04379_ ) );
BUF_X1 \mreg/_12736_ ( .A(\mreg/rf[21][29] ), .Z(\mreg/_04347_ ) );
BUF_X1 \mreg/_12737_ ( .A(\mreg/rf[20][29] ), .Z(\mreg/_04315_ ) );
BUF_X1 \mreg/_12738_ ( .A(\mreg/rf[19][29] ), .Z(\mreg/_04251_ ) );
BUF_X1 \mreg/_12739_ ( .A(\mreg/rf[18][29] ), .Z(\mreg/_04219_ ) );
BUF_X1 \mreg/_12740_ ( .A(\mreg/rf[17][29] ), .Z(\mreg/_04187_ ) );
BUF_X1 \mreg/_12741_ ( .A(\mreg/rf[16][29] ), .Z(\mreg/_04155_ ) );
BUF_X1 \mreg/_12742_ ( .A(\mreg/rf[15][29] ), .Z(\mreg/_04123_ ) );
BUF_X1 \mreg/_12743_ ( .A(\mreg/rf[14][29] ), .Z(\mreg/_04091_ ) );
BUF_X1 \mreg/_12744_ ( .A(\mreg/rf[13][29] ), .Z(\mreg/_04059_ ) );
BUF_X1 \mreg/_12745_ ( .A(\mreg/rf[12][29] ), .Z(\mreg/_04027_ ) );
BUF_X1 \mreg/_12746_ ( .A(\mreg/rf[11][29] ), .Z(\mreg/_03995_ ) );
BUF_X1 \mreg/_12747_ ( .A(\mreg/rf[10][29] ), .Z(\mreg/_03963_ ) );
BUF_X1 \mreg/_12748_ ( .A(\mreg/rf[9][29] ), .Z(\mreg/_04923_ ) );
BUF_X1 \mreg/_12749_ ( .A(\mreg/rf[8][29] ), .Z(\mreg/_04891_ ) );
BUF_X1 \mreg/_12750_ ( .A(\mreg/rf[7][29] ), .Z(\mreg/_04859_ ) );
BUF_X1 \mreg/_12751_ ( .A(\mreg/rf[6][29] ), .Z(\mreg/_04827_ ) );
BUF_X1 \mreg/_12752_ ( .A(\mreg/rf[5][29] ), .Z(\mreg/_04795_ ) );
BUF_X1 \mreg/_12753_ ( .A(\mreg/rf[4][29] ), .Z(\mreg/_04763_ ) );
BUF_X1 \mreg/_12754_ ( .A(\mreg/rf[3][29] ), .Z(\mreg/_04731_ ) );
BUF_X1 \mreg/_12755_ ( .A(\mreg/rf[2][29] ), .Z(\mreg/_04635_ ) );
BUF_X1 \mreg/_12756_ ( .A(\mreg/rf[1][29] ), .Z(\mreg/_04283_ ) );
BUF_X1 \mreg/_12757_ ( .A(\mreg/_03931_ ), .Z(\mem_wdata[29] ) );
BUF_X1 \mreg/_12758_ ( .A(\mreg/_00029_ ), .Z(\mreg/_00060_ ) );
BUF_X1 \mreg/_12759_ ( .A(\mreg/rf[30][30] ), .Z(\mreg/_04669_ ) );
BUF_X1 \mreg/_12760_ ( .A(\mreg/rf[29][30] ), .Z(\mreg/_04605_ ) );
BUF_X1 \mreg/_12761_ ( .A(\mreg/rf[28][30] ), .Z(\mreg/_04573_ ) );
BUF_X1 \mreg/_12762_ ( .A(\mreg/rf[27][30] ), .Z(\mreg/_04541_ ) );
BUF_X1 \mreg/_12763_ ( .A(\mreg/rf[26][30] ), .Z(\mreg/_04509_ ) );
BUF_X1 \mreg/_12764_ ( .A(\mreg/rf[25][30] ), .Z(\mreg/_04477_ ) );
BUF_X1 \mreg/_12765_ ( .A(\mreg/rf[24][30] ), .Z(\mreg/_04445_ ) );
BUF_X1 \mreg/_12766_ ( .A(\mreg/rf[23][30] ), .Z(\mreg/_04413_ ) );
BUF_X1 \mreg/_12767_ ( .A(\mreg/rf[22][30] ), .Z(\mreg/_04381_ ) );
BUF_X1 \mreg/_12768_ ( .A(\mreg/rf[21][30] ), .Z(\mreg/_04349_ ) );
BUF_X1 \mreg/_12769_ ( .A(\mreg/rf[20][30] ), .Z(\mreg/_04317_ ) );
BUF_X1 \mreg/_12770_ ( .A(\mreg/rf[19][30] ), .Z(\mreg/_04253_ ) );
BUF_X1 \mreg/_12771_ ( .A(\mreg/rf[18][30] ), .Z(\mreg/_04221_ ) );
BUF_X1 \mreg/_12772_ ( .A(\mreg/rf[17][30] ), .Z(\mreg/_04189_ ) );
BUF_X1 \mreg/_12773_ ( .A(\mreg/rf[16][30] ), .Z(\mreg/_04157_ ) );
BUF_X1 \mreg/_12774_ ( .A(\mreg/rf[15][30] ), .Z(\mreg/_04125_ ) );
BUF_X1 \mreg/_12775_ ( .A(\mreg/rf[14][30] ), .Z(\mreg/_04093_ ) );
BUF_X1 \mreg/_12776_ ( .A(\mreg/rf[13][30] ), .Z(\mreg/_04061_ ) );
BUF_X1 \mreg/_12777_ ( .A(\mreg/rf[12][30] ), .Z(\mreg/_04029_ ) );
BUF_X1 \mreg/_12778_ ( .A(\mreg/rf[11][30] ), .Z(\mreg/_03997_ ) );
BUF_X1 \mreg/_12779_ ( .A(\mreg/rf[10][30] ), .Z(\mreg/_03965_ ) );
BUF_X1 \mreg/_12780_ ( .A(\mreg/rf[9][30] ), .Z(\mreg/_04925_ ) );
BUF_X1 \mreg/_12781_ ( .A(\mreg/rf[8][30] ), .Z(\mreg/_04893_ ) );
BUF_X1 \mreg/_12782_ ( .A(\mreg/rf[7][30] ), .Z(\mreg/_04861_ ) );
BUF_X1 \mreg/_12783_ ( .A(\mreg/rf[6][30] ), .Z(\mreg/_04829_ ) );
BUF_X1 \mreg/_12784_ ( .A(\mreg/rf[5][30] ), .Z(\mreg/_04797_ ) );
BUF_X1 \mreg/_12785_ ( .A(\mreg/rf[4][30] ), .Z(\mreg/_04765_ ) );
BUF_X1 \mreg/_12786_ ( .A(\mreg/rf[3][30] ), .Z(\mreg/_04733_ ) );
BUF_X1 \mreg/_12787_ ( .A(\mreg/rf[2][30] ), .Z(\mreg/_04637_ ) );
BUF_X1 \mreg/_12788_ ( .A(\mreg/rf[1][30] ), .Z(\mreg/_04285_ ) );
BUF_X1 \mreg/_12789_ ( .A(\mreg/_03933_ ), .Z(\mem_wdata[30] ) );
BUF_X1 \mreg/_12790_ ( .A(\mreg/_00030_ ), .Z(\mreg/_00061_ ) );
BUF_X1 \mreg/_12791_ ( .A(\mreg/rf[30][31] ), .Z(\mreg/_04670_ ) );
BUF_X1 \mreg/_12792_ ( .A(\mreg/rf[29][31] ), .Z(\mreg/_04606_ ) );
BUF_X1 \mreg/_12793_ ( .A(\mreg/rf[28][31] ), .Z(\mreg/_04574_ ) );
BUF_X1 \mreg/_12794_ ( .A(\mreg/rf[27][31] ), .Z(\mreg/_04542_ ) );
BUF_X1 \mreg/_12795_ ( .A(\mreg/rf[26][31] ), .Z(\mreg/_04510_ ) );
BUF_X1 \mreg/_12796_ ( .A(\mreg/rf[25][31] ), .Z(\mreg/_04478_ ) );
BUF_X1 \mreg/_12797_ ( .A(\mreg/rf[24][31] ), .Z(\mreg/_04446_ ) );
BUF_X1 \mreg/_12798_ ( .A(\mreg/rf[23][31] ), .Z(\mreg/_04414_ ) );
BUF_X1 \mreg/_12799_ ( .A(\mreg/rf[22][31] ), .Z(\mreg/_04382_ ) );
BUF_X1 \mreg/_12800_ ( .A(\mreg/rf[21][31] ), .Z(\mreg/_04350_ ) );
BUF_X1 \mreg/_12801_ ( .A(\mreg/rf[20][31] ), .Z(\mreg/_04318_ ) );
BUF_X1 \mreg/_12802_ ( .A(\mreg/rf[19][31] ), .Z(\mreg/_04254_ ) );
BUF_X1 \mreg/_12803_ ( .A(\mreg/rf[18][31] ), .Z(\mreg/_04222_ ) );
BUF_X1 \mreg/_12804_ ( .A(\mreg/rf[17][31] ), .Z(\mreg/_04190_ ) );
BUF_X1 \mreg/_12805_ ( .A(\mreg/rf[16][31] ), .Z(\mreg/_04158_ ) );
BUF_X1 \mreg/_12806_ ( .A(\mreg/rf[15][31] ), .Z(\mreg/_04126_ ) );
BUF_X1 \mreg/_12807_ ( .A(\mreg/rf[14][31] ), .Z(\mreg/_04094_ ) );
BUF_X1 \mreg/_12808_ ( .A(\mreg/rf[13][31] ), .Z(\mreg/_04062_ ) );
BUF_X1 \mreg/_12809_ ( .A(\mreg/rf[12][31] ), .Z(\mreg/_04030_ ) );
BUF_X1 \mreg/_12810_ ( .A(\mreg/rf[11][31] ), .Z(\mreg/_03998_ ) );
BUF_X1 \mreg/_12811_ ( .A(\mreg/rf[10][31] ), .Z(\mreg/_03966_ ) );
BUF_X1 \mreg/_12812_ ( .A(\mreg/rf[9][31] ), .Z(\mreg/_04926_ ) );
BUF_X1 \mreg/_12813_ ( .A(\mreg/rf[8][31] ), .Z(\mreg/_04894_ ) );
BUF_X1 \mreg/_12814_ ( .A(\mreg/rf[7][31] ), .Z(\mreg/_04862_ ) );
BUF_X1 \mreg/_12815_ ( .A(\mreg/rf[6][31] ), .Z(\mreg/_04830_ ) );
BUF_X1 \mreg/_12816_ ( .A(\mreg/rf[5][31] ), .Z(\mreg/_04798_ ) );
BUF_X1 \mreg/_12817_ ( .A(\mreg/rf[4][31] ), .Z(\mreg/_04766_ ) );
BUF_X1 \mreg/_12818_ ( .A(\mreg/rf[3][31] ), .Z(\mreg/_04734_ ) );
BUF_X1 \mreg/_12819_ ( .A(\mreg/rf[2][31] ), .Z(\mreg/_04638_ ) );
BUF_X1 \mreg/_12820_ ( .A(\mreg/rf[1][31] ), .Z(\mreg/_04286_ ) );
BUF_X1 \mreg/_12821_ ( .A(\mreg/_03934_ ), .Z(\mem_wdata[31] ) );
BUF_X1 \mreg/_12822_ ( .A(\rs1[4] ), .Z(\mreg/_03872_ ) );
BUF_X1 \mreg/_12823_ ( .A(\rs1[1] ), .Z(\mreg/_03869_ ) );
BUF_X1 \mreg/_12824_ ( .A(\rs1[0] ), .Z(\mreg/_03868_ ) );
BUF_X1 \mreg/_12825_ ( .A(\rs1[3] ), .Z(\mreg/_03871_ ) );
BUF_X1 \mreg/_12826_ ( .A(\rs1[2] ), .Z(\mreg/_03870_ ) );
BUF_X1 \mreg/_12827_ ( .A(\mreg/_03878_ ), .Z(\src1[0] ) );
BUF_X1 \mreg/_12828_ ( .A(\mreg/_03889_ ), .Z(\src1[1] ) );
BUF_X1 \mreg/_12829_ ( .A(\mreg/_03900_ ), .Z(\src1[2] ) );
BUF_X1 \mreg/_12830_ ( .A(\mreg/_03903_ ), .Z(\src1[3] ) );
BUF_X1 \mreg/_12831_ ( .A(\mreg/_03904_ ), .Z(\src1[4] ) );
BUF_X1 \mreg/_12832_ ( .A(\mreg/_03905_ ), .Z(\src1[5] ) );
BUF_X1 \mreg/_12833_ ( .A(\mreg/_03906_ ), .Z(\src1[6] ) );
BUF_X1 \mreg/_12834_ ( .A(\mreg/_03907_ ), .Z(\src1[7] ) );
BUF_X1 \mreg/_12835_ ( .A(\mreg/_03908_ ), .Z(\src1[8] ) );
BUF_X1 \mreg/_12836_ ( .A(\mreg/_03909_ ), .Z(\src1[9] ) );
BUF_X1 \mreg/_12837_ ( .A(\mreg/_03879_ ), .Z(\src1[10] ) );
BUF_X1 \mreg/_12838_ ( .A(\mreg/_03880_ ), .Z(\src1[11] ) );
BUF_X1 \mreg/_12839_ ( .A(\mreg/_03881_ ), .Z(\src1[12] ) );
BUF_X1 \mreg/_12840_ ( .A(\mreg/_03882_ ), .Z(\src1[13] ) );
BUF_X1 \mreg/_12841_ ( .A(\mreg/_03883_ ), .Z(\src1[14] ) );
BUF_X1 \mreg/_12842_ ( .A(\mreg/_03884_ ), .Z(\src1[15] ) );
BUF_X1 \mreg/_12843_ ( .A(\mreg/_03885_ ), .Z(\src1[16] ) );
BUF_X1 \mreg/_12844_ ( .A(\mreg/_03886_ ), .Z(\src1[17] ) );
BUF_X1 \mreg/_12845_ ( .A(\mreg/_03887_ ), .Z(\src1[18] ) );
BUF_X1 \mreg/_12846_ ( .A(\mreg/_03888_ ), .Z(\src1[19] ) );
BUF_X1 \mreg/_12847_ ( .A(\mreg/_03890_ ), .Z(\src1[20] ) );
BUF_X1 \mreg/_12848_ ( .A(\mreg/_03891_ ), .Z(\src1[21] ) );
BUF_X1 \mreg/_12849_ ( .A(\mreg/_03892_ ), .Z(\src1[22] ) );
BUF_X1 \mreg/_12850_ ( .A(\mreg/_03893_ ), .Z(\src1[23] ) );
BUF_X1 \mreg/_12851_ ( .A(\mreg/_03894_ ), .Z(\src1[24] ) );
BUF_X1 \mreg/_12852_ ( .A(\mreg/_03895_ ), .Z(\src1[25] ) );
BUF_X1 \mreg/_12853_ ( .A(\mreg/_03896_ ), .Z(\src1[26] ) );
BUF_X1 \mreg/_12854_ ( .A(\mreg/_03897_ ), .Z(\src1[27] ) );
BUF_X1 \mreg/_12855_ ( .A(\mreg/_03898_ ), .Z(\src1[28] ) );
BUF_X1 \mreg/_12856_ ( .A(\mreg/_03899_ ), .Z(\src1[29] ) );
BUF_X1 \mreg/_12857_ ( .A(\mreg/_03901_ ), .Z(\src1[30] ) );
BUF_X1 \mreg/_12858_ ( .A(\mreg/_03902_ ), .Z(\src1[31] ) );
BUF_X1 \mreg/_12859_ ( .A(\result[0] ), .Z(\mreg/_04939_ ) );
BUF_X1 \mreg/_12860_ ( .A(\mreg/_00062_ ), .Z(\mreg/_05933_ ) );
BUF_X1 \mreg/_12861_ ( .A(\mreg/rf[31][1] ), .Z(\mreg/_04689_ ) );
BUF_X1 \mreg/_12862_ ( .A(\result[1] ), .Z(\mreg/_04950_ ) );
BUF_X1 \mreg/_12863_ ( .A(\mreg/_00063_ ), .Z(\mreg/_05934_ ) );
BUF_X1 \mreg/_12864_ ( .A(\mreg/rf[31][2] ), .Z(\mreg/_04700_ ) );
BUF_X1 \mreg/_12865_ ( .A(\result[2] ), .Z(\mreg/_04961_ ) );
BUF_X1 \mreg/_12866_ ( .A(\mreg/_00064_ ), .Z(\mreg/_05935_ ) );
BUF_X1 \mreg/_12867_ ( .A(\mreg/rf[31][3] ), .Z(\mreg/_04703_ ) );
BUF_X1 \mreg/_12868_ ( .A(\result[3] ), .Z(\mreg/_04964_ ) );
BUF_X1 \mreg/_12869_ ( .A(\mreg/_00065_ ), .Z(\mreg/_05936_ ) );
BUF_X1 \mreg/_12870_ ( .A(\mreg/rf[31][4] ), .Z(\mreg/_04704_ ) );
BUF_X1 \mreg/_12871_ ( .A(\result[4] ), .Z(\mreg/_04965_ ) );
BUF_X1 \mreg/_12872_ ( .A(\mreg/_00066_ ), .Z(\mreg/_05937_ ) );
BUF_X1 \mreg/_12873_ ( .A(\mreg/rf[31][5] ), .Z(\mreg/_04705_ ) );
BUF_X1 \mreg/_12874_ ( .A(\result[5] ), .Z(\mreg/_04966_ ) );
BUF_X1 \mreg/_12875_ ( .A(\mreg/_00067_ ), .Z(\mreg/_05938_ ) );
BUF_X1 \mreg/_12876_ ( .A(\mreg/rf[31][6] ), .Z(\mreg/_04706_ ) );
BUF_X1 \mreg/_12877_ ( .A(\result[6] ), .Z(\mreg/_04967_ ) );
BUF_X1 \mreg/_12878_ ( .A(\mreg/_00068_ ), .Z(\mreg/_05939_ ) );
BUF_X1 \mreg/_12879_ ( .A(\mreg/rf[31][7] ), .Z(\mreg/_04707_ ) );
BUF_X1 \mreg/_12880_ ( .A(\result[7] ), .Z(\mreg/_04968_ ) );
BUF_X1 \mreg/_12881_ ( .A(\mreg/_00069_ ), .Z(\mreg/_05940_ ) );
BUF_X1 \mreg/_12882_ ( .A(\mreg/rf[31][8] ), .Z(\mreg/_04708_ ) );
BUF_X1 \mreg/_12883_ ( .A(\result[8] ), .Z(\mreg/_04969_ ) );
BUF_X1 \mreg/_12884_ ( .A(\mreg/_00070_ ), .Z(\mreg/_05941_ ) );
BUF_X1 \mreg/_12885_ ( .A(\mreg/rf[31][9] ), .Z(\mreg/_04709_ ) );
BUF_X1 \mreg/_12886_ ( .A(\result[9] ), .Z(\mreg/_04970_ ) );
BUF_X1 \mreg/_12887_ ( .A(\mreg/_00071_ ), .Z(\mreg/_05942_ ) );
BUF_X1 \mreg/_12888_ ( .A(\mreg/rf[31][10] ), .Z(\mreg/_04679_ ) );
BUF_X1 \mreg/_12889_ ( .A(\result[10] ), .Z(\mreg/_04940_ ) );
BUF_X1 \mreg/_12890_ ( .A(\mreg/_00072_ ), .Z(\mreg/_05943_ ) );
BUF_X1 \mreg/_12891_ ( .A(\mreg/rf[31][11] ), .Z(\mreg/_04680_ ) );
BUF_X1 \mreg/_12892_ ( .A(\result[11] ), .Z(\mreg/_04941_ ) );
BUF_X1 \mreg/_12893_ ( .A(\mreg/_00073_ ), .Z(\mreg/_05944_ ) );
BUF_X1 \mreg/_12894_ ( .A(\mreg/rf[31][12] ), .Z(\mreg/_04681_ ) );
BUF_X1 \mreg/_12895_ ( .A(\result[12] ), .Z(\mreg/_04942_ ) );
BUF_X1 \mreg/_12896_ ( .A(\mreg/_00074_ ), .Z(\mreg/_05945_ ) );
BUF_X1 \mreg/_12897_ ( .A(\mreg/rf[31][13] ), .Z(\mreg/_04682_ ) );
BUF_X1 \mreg/_12898_ ( .A(\result[13] ), .Z(\mreg/_04943_ ) );
BUF_X1 \mreg/_12899_ ( .A(\mreg/_00075_ ), .Z(\mreg/_05946_ ) );
BUF_X1 \mreg/_12900_ ( .A(\mreg/rf[31][14] ), .Z(\mreg/_04683_ ) );
BUF_X1 \mreg/_12901_ ( .A(\result[14] ), .Z(\mreg/_04944_ ) );
BUF_X1 \mreg/_12902_ ( .A(\mreg/_00076_ ), .Z(\mreg/_05947_ ) );
BUF_X1 \mreg/_12903_ ( .A(\mreg/rf[31][15] ), .Z(\mreg/_04684_ ) );
BUF_X1 \mreg/_12904_ ( .A(\result[15] ), .Z(\mreg/_04945_ ) );
BUF_X1 \mreg/_12905_ ( .A(\mreg/_00077_ ), .Z(\mreg/_05948_ ) );
BUF_X1 \mreg/_12906_ ( .A(\mreg/rf[31][16] ), .Z(\mreg/_04685_ ) );
BUF_X1 \mreg/_12907_ ( .A(\result[16] ), .Z(\mreg/_04946_ ) );
BUF_X1 \mreg/_12908_ ( .A(\mreg/_00078_ ), .Z(\mreg/_05949_ ) );
BUF_X1 \mreg/_12909_ ( .A(\mreg/rf[31][17] ), .Z(\mreg/_04686_ ) );
BUF_X1 \mreg/_12910_ ( .A(\result[17] ), .Z(\mreg/_04947_ ) );
BUF_X1 \mreg/_12911_ ( .A(\mreg/_00079_ ), .Z(\mreg/_05950_ ) );
BUF_X1 \mreg/_12912_ ( .A(\mreg/rf[31][18] ), .Z(\mreg/_04687_ ) );
BUF_X1 \mreg/_12913_ ( .A(\result[18] ), .Z(\mreg/_04948_ ) );
BUF_X1 \mreg/_12914_ ( .A(\mreg/_00080_ ), .Z(\mreg/_05951_ ) );
BUF_X1 \mreg/_12915_ ( .A(\mreg/rf[31][19] ), .Z(\mreg/_04688_ ) );
BUF_X1 \mreg/_12916_ ( .A(\result[19] ), .Z(\mreg/_04949_ ) );
BUF_X1 \mreg/_12917_ ( .A(\mreg/_00081_ ), .Z(\mreg/_05952_ ) );
BUF_X1 \mreg/_12918_ ( .A(\mreg/rf[31][20] ), .Z(\mreg/_04690_ ) );
BUF_X1 \mreg/_12919_ ( .A(\result[20] ), .Z(\mreg/_04951_ ) );
BUF_X1 \mreg/_12920_ ( .A(\mreg/_00082_ ), .Z(\mreg/_05953_ ) );
BUF_X1 \mreg/_12921_ ( .A(\mreg/rf[31][21] ), .Z(\mreg/_04691_ ) );
BUF_X1 \mreg/_12922_ ( .A(\result[21] ), .Z(\mreg/_04952_ ) );
BUF_X1 \mreg/_12923_ ( .A(\mreg/_00083_ ), .Z(\mreg/_05954_ ) );
BUF_X1 \mreg/_12924_ ( .A(\mreg/rf[31][22] ), .Z(\mreg/_04692_ ) );
BUF_X1 \mreg/_12925_ ( .A(\result[22] ), .Z(\mreg/_04953_ ) );
BUF_X1 \mreg/_12926_ ( .A(\mreg/_00084_ ), .Z(\mreg/_05955_ ) );
BUF_X1 \mreg/_12927_ ( .A(\mreg/rf[31][23] ), .Z(\mreg/_04693_ ) );
BUF_X1 \mreg/_12928_ ( .A(\result[23] ), .Z(\mreg/_04954_ ) );
BUF_X1 \mreg/_12929_ ( .A(\mreg/_00085_ ), .Z(\mreg/_05956_ ) );
BUF_X1 \mreg/_12930_ ( .A(\mreg/rf[31][24] ), .Z(\mreg/_04694_ ) );
BUF_X1 \mreg/_12931_ ( .A(\result[24] ), .Z(\mreg/_04955_ ) );
BUF_X1 \mreg/_12932_ ( .A(\mreg/_00086_ ), .Z(\mreg/_05957_ ) );
BUF_X1 \mreg/_12933_ ( .A(\mreg/rf[31][25] ), .Z(\mreg/_04695_ ) );
BUF_X1 \mreg/_12934_ ( .A(\result[25] ), .Z(\mreg/_04956_ ) );
BUF_X1 \mreg/_12935_ ( .A(\mreg/_00087_ ), .Z(\mreg/_05958_ ) );
BUF_X1 \mreg/_12936_ ( .A(\mreg/rf[31][26] ), .Z(\mreg/_04696_ ) );
BUF_X1 \mreg/_12937_ ( .A(\result[26] ), .Z(\mreg/_04957_ ) );
BUF_X1 \mreg/_12938_ ( .A(\mreg/_00088_ ), .Z(\mreg/_05959_ ) );
BUF_X1 \mreg/_12939_ ( .A(\mreg/rf[31][27] ), .Z(\mreg/_04697_ ) );
BUF_X1 \mreg/_12940_ ( .A(\result[27] ), .Z(\mreg/_04958_ ) );
BUF_X1 \mreg/_12941_ ( .A(\mreg/_00089_ ), .Z(\mreg/_05960_ ) );
BUF_X1 \mreg/_12942_ ( .A(\mreg/rf[31][28] ), .Z(\mreg/_04698_ ) );
BUF_X1 \mreg/_12943_ ( .A(\result[28] ), .Z(\mreg/_04959_ ) );
BUF_X1 \mreg/_12944_ ( .A(\mreg/_00090_ ), .Z(\mreg/_05961_ ) );
BUF_X1 \mreg/_12945_ ( .A(\mreg/rf[31][29] ), .Z(\mreg/_04699_ ) );
BUF_X1 \mreg/_12946_ ( .A(\result[29] ), .Z(\mreg/_04960_ ) );
BUF_X1 \mreg/_12947_ ( .A(\mreg/_00091_ ), .Z(\mreg/_05962_ ) );
BUF_X1 \mreg/_12948_ ( .A(\mreg/rf[31][30] ), .Z(\mreg/_04701_ ) );
BUF_X1 \mreg/_12949_ ( .A(\result[30] ), .Z(\mreg/_04962_ ) );
BUF_X1 \mreg/_12950_ ( .A(\mreg/_00092_ ), .Z(\mreg/_05963_ ) );
BUF_X1 \mreg/_12951_ ( .A(\mreg/rf[31][31] ), .Z(\mreg/_04702_ ) );
BUF_X1 \mreg/_12952_ ( .A(\result[31] ), .Z(\mreg/_04963_ ) );
BUF_X1 \mreg/_12953_ ( .A(\mreg/_00093_ ), .Z(\mreg/_05964_ ) );
BUF_X1 \mreg/_12954_ ( .A(\mreg/_00094_ ), .Z(\mreg/_05965_ ) );
BUF_X1 \mreg/_12955_ ( .A(\mreg/_00095_ ), .Z(\mreg/_05966_ ) );
BUF_X1 \mreg/_12956_ ( .A(\mreg/_00096_ ), .Z(\mreg/_05967_ ) );
BUF_X1 \mreg/_12957_ ( .A(\mreg/_00097_ ), .Z(\mreg/_05968_ ) );
BUF_X1 \mreg/_12958_ ( .A(\mreg/_00098_ ), .Z(\mreg/_05969_ ) );
BUF_X1 \mreg/_12959_ ( .A(\mreg/_00099_ ), .Z(\mreg/_05970_ ) );
BUF_X1 \mreg/_12960_ ( .A(\mreg/_00100_ ), .Z(\mreg/_05971_ ) );
BUF_X1 \mreg/_12961_ ( .A(\mreg/_00101_ ), .Z(\mreg/_05972_ ) );
BUF_X1 \mreg/_12962_ ( .A(\mreg/_00102_ ), .Z(\mreg/_05973_ ) );
BUF_X1 \mreg/_12963_ ( .A(\mreg/_00103_ ), .Z(\mreg/_05974_ ) );
BUF_X1 \mreg/_12964_ ( .A(\mreg/_00104_ ), .Z(\mreg/_05975_ ) );
BUF_X1 \mreg/_12965_ ( .A(\mreg/_00105_ ), .Z(\mreg/_05976_ ) );
BUF_X1 \mreg/_12966_ ( .A(\mreg/_00106_ ), .Z(\mreg/_05977_ ) );
BUF_X1 \mreg/_12967_ ( .A(\mreg/_00107_ ), .Z(\mreg/_05978_ ) );
BUF_X1 \mreg/_12968_ ( .A(\mreg/_00108_ ), .Z(\mreg/_05979_ ) );
BUF_X1 \mreg/_12969_ ( .A(\mreg/_00109_ ), .Z(\mreg/_05980_ ) );
BUF_X1 \mreg/_12970_ ( .A(\mreg/_00110_ ), .Z(\mreg/_05981_ ) );
BUF_X1 \mreg/_12971_ ( .A(\mreg/_00111_ ), .Z(\mreg/_05982_ ) );
BUF_X1 \mreg/_12972_ ( .A(\mreg/_00112_ ), .Z(\mreg/_05983_ ) );
BUF_X1 \mreg/_12973_ ( .A(\mreg/_00113_ ), .Z(\mreg/_05984_ ) );
BUF_X1 \mreg/_12974_ ( .A(\mreg/_00114_ ), .Z(\mreg/_05985_ ) );
BUF_X1 \mreg/_12975_ ( .A(\mreg/_00115_ ), .Z(\mreg/_05986_ ) );
BUF_X1 \mreg/_12976_ ( .A(\mreg/_00116_ ), .Z(\mreg/_05987_ ) );
BUF_X1 \mreg/_12977_ ( .A(\mreg/_00117_ ), .Z(\mreg/_05988_ ) );
BUF_X1 \mreg/_12978_ ( .A(\mreg/_00118_ ), .Z(\mreg/_05989_ ) );
BUF_X1 \mreg/_12979_ ( .A(\mreg/_00119_ ), .Z(\mreg/_05990_ ) );
BUF_X1 \mreg/_12980_ ( .A(\mreg/_00120_ ), .Z(\mreg/_05991_ ) );
BUF_X1 \mreg/_12981_ ( .A(\mreg/_00121_ ), .Z(\mreg/_05992_ ) );
BUF_X1 \mreg/_12982_ ( .A(\mreg/_00122_ ), .Z(\mreg/_05993_ ) );
BUF_X1 \mreg/_12983_ ( .A(\mreg/_00123_ ), .Z(\mreg/_05994_ ) );
BUF_X1 \mreg/_12984_ ( .A(\mreg/_00124_ ), .Z(\mreg/_05995_ ) );
BUF_X1 \mreg/_12985_ ( .A(\mreg/_00125_ ), .Z(\mreg/_05996_ ) );
BUF_X1 \mreg/_12986_ ( .A(\mreg/_00126_ ), .Z(\mreg/_05997_ ) );
BUF_X1 \mreg/_12987_ ( .A(\mreg/_00127_ ), .Z(\mreg/_05998_ ) );
BUF_X1 \mreg/_12988_ ( .A(\mreg/_00128_ ), .Z(\mreg/_05999_ ) );
BUF_X1 \mreg/_12989_ ( .A(\mreg/_00129_ ), .Z(\mreg/_06000_ ) );
BUF_X1 \mreg/_12990_ ( .A(\mreg/_00130_ ), .Z(\mreg/_06001_ ) );
BUF_X1 \mreg/_12991_ ( .A(\mreg/_00131_ ), .Z(\mreg/_06002_ ) );
BUF_X1 \mreg/_12992_ ( .A(\mreg/_00132_ ), .Z(\mreg/_06003_ ) );
BUF_X1 \mreg/_12993_ ( .A(\mreg/_00133_ ), .Z(\mreg/_06004_ ) );
BUF_X1 \mreg/_12994_ ( .A(\mreg/_00134_ ), .Z(\mreg/_06005_ ) );
BUF_X1 \mreg/_12995_ ( .A(\mreg/_00135_ ), .Z(\mreg/_06006_ ) );
BUF_X1 \mreg/_12996_ ( .A(\mreg/_00136_ ), .Z(\mreg/_06007_ ) );
BUF_X1 \mreg/_12997_ ( .A(\mreg/_00137_ ), .Z(\mreg/_06008_ ) );
BUF_X1 \mreg/_12998_ ( .A(\mreg/_00138_ ), .Z(\mreg/_06009_ ) );
BUF_X1 \mreg/_12999_ ( .A(\mreg/_00139_ ), .Z(\mreg/_06010_ ) );
BUF_X1 \mreg/_13000_ ( .A(\mreg/_00140_ ), .Z(\mreg/_06011_ ) );
BUF_X1 \mreg/_13001_ ( .A(\mreg/_00141_ ), .Z(\mreg/_06012_ ) );
BUF_X1 \mreg/_13002_ ( .A(\mreg/_00142_ ), .Z(\mreg/_06013_ ) );
BUF_X1 \mreg/_13003_ ( .A(\mreg/_00143_ ), .Z(\mreg/_06014_ ) );
BUF_X1 \mreg/_13004_ ( .A(\mreg/_00144_ ), .Z(\mreg/_06015_ ) );
BUF_X1 \mreg/_13005_ ( .A(\mreg/_00145_ ), .Z(\mreg/_06016_ ) );
BUF_X1 \mreg/_13006_ ( .A(\mreg/_00146_ ), .Z(\mreg/_06017_ ) );
BUF_X1 \mreg/_13007_ ( .A(\mreg/_00147_ ), .Z(\mreg/_06018_ ) );
BUF_X1 \mreg/_13008_ ( .A(\mreg/_00148_ ), .Z(\mreg/_06019_ ) );
BUF_X1 \mreg/_13009_ ( .A(\mreg/_00149_ ), .Z(\mreg/_06020_ ) );
BUF_X1 \mreg/_13010_ ( .A(\mreg/_00150_ ), .Z(\mreg/_06021_ ) );
BUF_X1 \mreg/_13011_ ( .A(\mreg/_00151_ ), .Z(\mreg/_06022_ ) );
BUF_X1 \mreg/_13012_ ( .A(\mreg/_00152_ ), .Z(\mreg/_06023_ ) );
BUF_X1 \mreg/_13013_ ( .A(\mreg/_00153_ ), .Z(\mreg/_06024_ ) );
BUF_X1 \mreg/_13014_ ( .A(\mreg/_00154_ ), .Z(\mreg/_06025_ ) );
BUF_X1 \mreg/_13015_ ( .A(\mreg/_00155_ ), .Z(\mreg/_06026_ ) );
BUF_X1 \mreg/_13016_ ( .A(\mreg/_00156_ ), .Z(\mreg/_06027_ ) );
BUF_X1 \mreg/_13017_ ( .A(\mreg/_00157_ ), .Z(\mreg/_06028_ ) );
BUF_X1 \mreg/_13018_ ( .A(\mreg/_00158_ ), .Z(\mreg/_06029_ ) );
BUF_X1 \mreg/_13019_ ( .A(\mreg/_00159_ ), .Z(\mreg/_06030_ ) );
BUF_X1 \mreg/_13020_ ( .A(\mreg/_00160_ ), .Z(\mreg/_06031_ ) );
BUF_X1 \mreg/_13021_ ( .A(\mreg/_00161_ ), .Z(\mreg/_06032_ ) );
BUF_X1 \mreg/_13022_ ( .A(\mreg/_00162_ ), .Z(\mreg/_06033_ ) );
BUF_X1 \mreg/_13023_ ( .A(\mreg/_00163_ ), .Z(\mreg/_06034_ ) );
BUF_X1 \mreg/_13024_ ( .A(\mreg/_00164_ ), .Z(\mreg/_06035_ ) );
BUF_X1 \mreg/_13025_ ( .A(\mreg/_00165_ ), .Z(\mreg/_06036_ ) );
BUF_X1 \mreg/_13026_ ( .A(\mreg/_00166_ ), .Z(\mreg/_06037_ ) );
BUF_X1 \mreg/_13027_ ( .A(\mreg/_00167_ ), .Z(\mreg/_06038_ ) );
BUF_X1 \mreg/_13028_ ( .A(\mreg/_00168_ ), .Z(\mreg/_06039_ ) );
BUF_X1 \mreg/_13029_ ( .A(\mreg/_00169_ ), .Z(\mreg/_06040_ ) );
BUF_X1 \mreg/_13030_ ( .A(\mreg/_00170_ ), .Z(\mreg/_06041_ ) );
BUF_X1 \mreg/_13031_ ( .A(\mreg/_00171_ ), .Z(\mreg/_06042_ ) );
BUF_X1 \mreg/_13032_ ( .A(\mreg/_00172_ ), .Z(\mreg/_06043_ ) );
BUF_X1 \mreg/_13033_ ( .A(\mreg/_00173_ ), .Z(\mreg/_06044_ ) );
BUF_X1 \mreg/_13034_ ( .A(\mreg/_00174_ ), .Z(\mreg/_06045_ ) );
BUF_X1 \mreg/_13035_ ( .A(\mreg/_00175_ ), .Z(\mreg/_06046_ ) );
BUF_X1 \mreg/_13036_ ( .A(\mreg/_00176_ ), .Z(\mreg/_06047_ ) );
BUF_X1 \mreg/_13037_ ( .A(\mreg/_00177_ ), .Z(\mreg/_06048_ ) );
BUF_X1 \mreg/_13038_ ( .A(\mreg/_00178_ ), .Z(\mreg/_06049_ ) );
BUF_X1 \mreg/_13039_ ( .A(\mreg/_00179_ ), .Z(\mreg/_06050_ ) );
BUF_X1 \mreg/_13040_ ( .A(\mreg/_00180_ ), .Z(\mreg/_06051_ ) );
BUF_X1 \mreg/_13041_ ( .A(\mreg/_00181_ ), .Z(\mreg/_06052_ ) );
BUF_X1 \mreg/_13042_ ( .A(\mreg/_00182_ ), .Z(\mreg/_06053_ ) );
BUF_X1 \mreg/_13043_ ( .A(\mreg/_00183_ ), .Z(\mreg/_06054_ ) );
BUF_X1 \mreg/_13044_ ( .A(\mreg/_00184_ ), .Z(\mreg/_06055_ ) );
BUF_X1 \mreg/_13045_ ( .A(\mreg/_00185_ ), .Z(\mreg/_06056_ ) );
BUF_X1 \mreg/_13046_ ( .A(\mreg/_00186_ ), .Z(\mreg/_06057_ ) );
BUF_X1 \mreg/_13047_ ( .A(\mreg/_00187_ ), .Z(\mreg/_06058_ ) );
BUF_X1 \mreg/_13048_ ( .A(\mreg/_00188_ ), .Z(\mreg/_06059_ ) );
BUF_X1 \mreg/_13049_ ( .A(\mreg/_00189_ ), .Z(\mreg/_06060_ ) );
BUF_X1 \mreg/_13050_ ( .A(\mreg/_00190_ ), .Z(\mreg/_06061_ ) );
BUF_X1 \mreg/_13051_ ( .A(\mreg/_00191_ ), .Z(\mreg/_06062_ ) );
BUF_X1 \mreg/_13052_ ( .A(\mreg/_00192_ ), .Z(\mreg/_06063_ ) );
BUF_X1 \mreg/_13053_ ( .A(\mreg/_00193_ ), .Z(\mreg/_06064_ ) );
BUF_X1 \mreg/_13054_ ( .A(\mreg/_00194_ ), .Z(\mreg/_06065_ ) );
BUF_X1 \mreg/_13055_ ( .A(\mreg/_00195_ ), .Z(\mreg/_06066_ ) );
BUF_X1 \mreg/_13056_ ( .A(\mreg/_00196_ ), .Z(\mreg/_06067_ ) );
BUF_X1 \mreg/_13057_ ( .A(\mreg/_00197_ ), .Z(\mreg/_06068_ ) );
BUF_X1 \mreg/_13058_ ( .A(\mreg/_00198_ ), .Z(\mreg/_06069_ ) );
BUF_X1 \mreg/_13059_ ( .A(\mreg/_00199_ ), .Z(\mreg/_06070_ ) );
BUF_X1 \mreg/_13060_ ( .A(\mreg/_00200_ ), .Z(\mreg/_06071_ ) );
BUF_X1 \mreg/_13061_ ( .A(\mreg/_00201_ ), .Z(\mreg/_06072_ ) );
BUF_X1 \mreg/_13062_ ( .A(\mreg/_00202_ ), .Z(\mreg/_06073_ ) );
BUF_X1 \mreg/_13063_ ( .A(\mreg/_00203_ ), .Z(\mreg/_06074_ ) );
BUF_X1 \mreg/_13064_ ( .A(\mreg/_00204_ ), .Z(\mreg/_06075_ ) );
BUF_X1 \mreg/_13065_ ( .A(\mreg/_00205_ ), .Z(\mreg/_06076_ ) );
BUF_X1 \mreg/_13066_ ( .A(\mreg/_00206_ ), .Z(\mreg/_06077_ ) );
BUF_X1 \mreg/_13067_ ( .A(\mreg/_00207_ ), .Z(\mreg/_06078_ ) );
BUF_X1 \mreg/_13068_ ( .A(\mreg/_00208_ ), .Z(\mreg/_06079_ ) );
BUF_X1 \mreg/_13069_ ( .A(\mreg/_00209_ ), .Z(\mreg/_06080_ ) );
BUF_X1 \mreg/_13070_ ( .A(\mreg/_00210_ ), .Z(\mreg/_06081_ ) );
BUF_X1 \mreg/_13071_ ( .A(\mreg/_00211_ ), .Z(\mreg/_06082_ ) );
BUF_X1 \mreg/_13072_ ( .A(\mreg/_00212_ ), .Z(\mreg/_06083_ ) );
BUF_X1 \mreg/_13073_ ( .A(\mreg/_00213_ ), .Z(\mreg/_06084_ ) );
BUF_X1 \mreg/_13074_ ( .A(\mreg/_00214_ ), .Z(\mreg/_06085_ ) );
BUF_X1 \mreg/_13075_ ( .A(\mreg/_00215_ ), .Z(\mreg/_06086_ ) );
BUF_X1 \mreg/_13076_ ( .A(\mreg/_00216_ ), .Z(\mreg/_06087_ ) );
BUF_X1 \mreg/_13077_ ( .A(\mreg/_00217_ ), .Z(\mreg/_06088_ ) );
BUF_X1 \mreg/_13078_ ( .A(\mreg/_00218_ ), .Z(\mreg/_06089_ ) );
BUF_X1 \mreg/_13079_ ( .A(\mreg/_00219_ ), .Z(\mreg/_06090_ ) );
BUF_X1 \mreg/_13080_ ( .A(\mreg/_00220_ ), .Z(\mreg/_06091_ ) );
BUF_X1 \mreg/_13081_ ( .A(\mreg/_00221_ ), .Z(\mreg/_06092_ ) );
BUF_X1 \mreg/_13082_ ( .A(\mreg/_00222_ ), .Z(\mreg/_06093_ ) );
BUF_X1 \mreg/_13083_ ( .A(\mreg/_00223_ ), .Z(\mreg/_06094_ ) );
BUF_X1 \mreg/_13084_ ( .A(\mreg/_00224_ ), .Z(\mreg/_06095_ ) );
BUF_X1 \mreg/_13085_ ( .A(\mreg/_00225_ ), .Z(\mreg/_06096_ ) );
BUF_X1 \mreg/_13086_ ( .A(\mreg/_00226_ ), .Z(\mreg/_06097_ ) );
BUF_X1 \mreg/_13087_ ( .A(\mreg/_00227_ ), .Z(\mreg/_06098_ ) );
BUF_X1 \mreg/_13088_ ( .A(\mreg/_00228_ ), .Z(\mreg/_06099_ ) );
BUF_X1 \mreg/_13089_ ( .A(\mreg/_00229_ ), .Z(\mreg/_06100_ ) );
BUF_X1 \mreg/_13090_ ( .A(\mreg/_00230_ ), .Z(\mreg/_06101_ ) );
BUF_X1 \mreg/_13091_ ( .A(\mreg/_00231_ ), .Z(\mreg/_06102_ ) );
BUF_X1 \mreg/_13092_ ( .A(\mreg/_00232_ ), .Z(\mreg/_06103_ ) );
BUF_X1 \mreg/_13093_ ( .A(\mreg/_00233_ ), .Z(\mreg/_06104_ ) );
BUF_X1 \mreg/_13094_ ( .A(\mreg/_00234_ ), .Z(\mreg/_06105_ ) );
BUF_X1 \mreg/_13095_ ( .A(\mreg/_00235_ ), .Z(\mreg/_06106_ ) );
BUF_X1 \mreg/_13096_ ( .A(\mreg/_00236_ ), .Z(\mreg/_06107_ ) );
BUF_X1 \mreg/_13097_ ( .A(\mreg/_00237_ ), .Z(\mreg/_06108_ ) );
BUF_X1 \mreg/_13098_ ( .A(\mreg/_00238_ ), .Z(\mreg/_06109_ ) );
BUF_X1 \mreg/_13099_ ( .A(\mreg/_00239_ ), .Z(\mreg/_06110_ ) );
BUF_X1 \mreg/_13100_ ( .A(\mreg/_00240_ ), .Z(\mreg/_06111_ ) );
BUF_X1 \mreg/_13101_ ( .A(\mreg/_00241_ ), .Z(\mreg/_06112_ ) );
BUF_X1 \mreg/_13102_ ( .A(\mreg/_00242_ ), .Z(\mreg/_06113_ ) );
BUF_X1 \mreg/_13103_ ( .A(\mreg/_00243_ ), .Z(\mreg/_06114_ ) );
BUF_X1 \mreg/_13104_ ( .A(\mreg/_00244_ ), .Z(\mreg/_06115_ ) );
BUF_X1 \mreg/_13105_ ( .A(\mreg/_00245_ ), .Z(\mreg/_06116_ ) );
BUF_X1 \mreg/_13106_ ( .A(\mreg/_00246_ ), .Z(\mreg/_06117_ ) );
BUF_X1 \mreg/_13107_ ( .A(\mreg/_00247_ ), .Z(\mreg/_06118_ ) );
BUF_X1 \mreg/_13108_ ( .A(\mreg/_00248_ ), .Z(\mreg/_06119_ ) );
BUF_X1 \mreg/_13109_ ( .A(\mreg/_00249_ ), .Z(\mreg/_06120_ ) );
BUF_X1 \mreg/_13110_ ( .A(\mreg/_00250_ ), .Z(\mreg/_06121_ ) );
BUF_X1 \mreg/_13111_ ( .A(\mreg/_00251_ ), .Z(\mreg/_06122_ ) );
BUF_X1 \mreg/_13112_ ( .A(\mreg/_00252_ ), .Z(\mreg/_06123_ ) );
BUF_X1 \mreg/_13113_ ( .A(\mreg/_00253_ ), .Z(\mreg/_06124_ ) );
BUF_X1 \mreg/_13114_ ( .A(\mreg/_00254_ ), .Z(\mreg/_06125_ ) );
BUF_X1 \mreg/_13115_ ( .A(\mreg/_00255_ ), .Z(\mreg/_06126_ ) );
BUF_X1 \mreg/_13116_ ( .A(\mreg/_00256_ ), .Z(\mreg/_06127_ ) );
BUF_X1 \mreg/_13117_ ( .A(\mreg/_00257_ ), .Z(\mreg/_06128_ ) );
BUF_X1 \mreg/_13118_ ( .A(\mreg/_00258_ ), .Z(\mreg/_06129_ ) );
BUF_X1 \mreg/_13119_ ( .A(\mreg/_00259_ ), .Z(\mreg/_06130_ ) );
BUF_X1 \mreg/_13120_ ( .A(\mreg/_00260_ ), .Z(\mreg/_06131_ ) );
BUF_X1 \mreg/_13121_ ( .A(\mreg/_00261_ ), .Z(\mreg/_06132_ ) );
BUF_X1 \mreg/_13122_ ( .A(\mreg/_00262_ ), .Z(\mreg/_06133_ ) );
BUF_X1 \mreg/_13123_ ( .A(\mreg/_00263_ ), .Z(\mreg/_06134_ ) );
BUF_X1 \mreg/_13124_ ( .A(\mreg/_00264_ ), .Z(\mreg/_06135_ ) );
BUF_X1 \mreg/_13125_ ( .A(\mreg/_00265_ ), .Z(\mreg/_06136_ ) );
BUF_X1 \mreg/_13126_ ( .A(\mreg/_00266_ ), .Z(\mreg/_06137_ ) );
BUF_X1 \mreg/_13127_ ( .A(\mreg/_00267_ ), .Z(\mreg/_06138_ ) );
BUF_X1 \mreg/_13128_ ( .A(\mreg/_00268_ ), .Z(\mreg/_06139_ ) );
BUF_X1 \mreg/_13129_ ( .A(\mreg/_00269_ ), .Z(\mreg/_06140_ ) );
BUF_X1 \mreg/_13130_ ( .A(\mreg/_00270_ ), .Z(\mreg/_06141_ ) );
BUF_X1 \mreg/_13131_ ( .A(\mreg/_00271_ ), .Z(\mreg/_06142_ ) );
BUF_X1 \mreg/_13132_ ( .A(\mreg/_00272_ ), .Z(\mreg/_06143_ ) );
BUF_X1 \mreg/_13133_ ( .A(\mreg/_00273_ ), .Z(\mreg/_06144_ ) );
BUF_X1 \mreg/_13134_ ( .A(\mreg/_00274_ ), .Z(\mreg/_06145_ ) );
BUF_X1 \mreg/_13135_ ( .A(\mreg/_00275_ ), .Z(\mreg/_06146_ ) );
BUF_X1 \mreg/_13136_ ( .A(\mreg/_00276_ ), .Z(\mreg/_06147_ ) );
BUF_X1 \mreg/_13137_ ( .A(\mreg/_00277_ ), .Z(\mreg/_06148_ ) );
BUF_X1 \mreg/_13138_ ( .A(\mreg/_00278_ ), .Z(\mreg/_06149_ ) );
BUF_X1 \mreg/_13139_ ( .A(\mreg/_00279_ ), .Z(\mreg/_06150_ ) );
BUF_X1 \mreg/_13140_ ( .A(\mreg/_00280_ ), .Z(\mreg/_06151_ ) );
BUF_X1 \mreg/_13141_ ( .A(\mreg/_00281_ ), .Z(\mreg/_06152_ ) );
BUF_X1 \mreg/_13142_ ( .A(\mreg/_00282_ ), .Z(\mreg/_06153_ ) );
BUF_X1 \mreg/_13143_ ( .A(\mreg/_00283_ ), .Z(\mreg/_06154_ ) );
BUF_X1 \mreg/_13144_ ( .A(\mreg/_00284_ ), .Z(\mreg/_06155_ ) );
BUF_X1 \mreg/_13145_ ( .A(\mreg/_00285_ ), .Z(\mreg/_06156_ ) );
BUF_X1 \mreg/_13146_ ( .A(\mreg/_00286_ ), .Z(\mreg/_06157_ ) );
BUF_X1 \mreg/_13147_ ( .A(\mreg/_00287_ ), .Z(\mreg/_06158_ ) );
BUF_X1 \mreg/_13148_ ( .A(\mreg/_00288_ ), .Z(\mreg/_06159_ ) );
BUF_X1 \mreg/_13149_ ( .A(\mreg/_00289_ ), .Z(\mreg/_06160_ ) );
BUF_X1 \mreg/_13150_ ( .A(\mreg/_00290_ ), .Z(\mreg/_06161_ ) );
BUF_X1 \mreg/_13151_ ( .A(\mreg/_00291_ ), .Z(\mreg/_06162_ ) );
BUF_X1 \mreg/_13152_ ( .A(\mreg/_00292_ ), .Z(\mreg/_06163_ ) );
BUF_X1 \mreg/_13153_ ( .A(\mreg/_00293_ ), .Z(\mreg/_06164_ ) );
BUF_X1 \mreg/_13154_ ( .A(\mreg/_00294_ ), .Z(\mreg/_06165_ ) );
BUF_X1 \mreg/_13155_ ( .A(\mreg/_00295_ ), .Z(\mreg/_06166_ ) );
BUF_X1 \mreg/_13156_ ( .A(\mreg/_00296_ ), .Z(\mreg/_06167_ ) );
BUF_X1 \mreg/_13157_ ( .A(\mreg/_00297_ ), .Z(\mreg/_06168_ ) );
BUF_X1 \mreg/_13158_ ( .A(\mreg/_00298_ ), .Z(\mreg/_06169_ ) );
BUF_X1 \mreg/_13159_ ( .A(\mreg/_00299_ ), .Z(\mreg/_06170_ ) );
BUF_X1 \mreg/_13160_ ( .A(\mreg/_00300_ ), .Z(\mreg/_06171_ ) );
BUF_X1 \mreg/_13161_ ( .A(\mreg/_00301_ ), .Z(\mreg/_06172_ ) );
BUF_X1 \mreg/_13162_ ( .A(\mreg/_00302_ ), .Z(\mreg/_06173_ ) );
BUF_X1 \mreg/_13163_ ( .A(\mreg/_00303_ ), .Z(\mreg/_06174_ ) );
BUF_X1 \mreg/_13164_ ( .A(\mreg/_00304_ ), .Z(\mreg/_06175_ ) );
BUF_X1 \mreg/_13165_ ( .A(\mreg/_00305_ ), .Z(\mreg/_06176_ ) );
BUF_X1 \mreg/_13166_ ( .A(\mreg/_00306_ ), .Z(\mreg/_06177_ ) );
BUF_X1 \mreg/_13167_ ( .A(\mreg/_00307_ ), .Z(\mreg/_06178_ ) );
BUF_X1 \mreg/_13168_ ( .A(\mreg/_00308_ ), .Z(\mreg/_06179_ ) );
BUF_X1 \mreg/_13169_ ( .A(\mreg/_00309_ ), .Z(\mreg/_06180_ ) );
BUF_X1 \mreg/_13170_ ( .A(\mreg/_00310_ ), .Z(\mreg/_06181_ ) );
BUF_X1 \mreg/_13171_ ( .A(\mreg/_00311_ ), .Z(\mreg/_06182_ ) );
BUF_X1 \mreg/_13172_ ( .A(\mreg/_00312_ ), .Z(\mreg/_06183_ ) );
BUF_X1 \mreg/_13173_ ( .A(\mreg/_00313_ ), .Z(\mreg/_06184_ ) );
BUF_X1 \mreg/_13174_ ( .A(\mreg/_00314_ ), .Z(\mreg/_06185_ ) );
BUF_X1 \mreg/_13175_ ( .A(\mreg/_00315_ ), .Z(\mreg/_06186_ ) );
BUF_X1 \mreg/_13176_ ( .A(\mreg/_00316_ ), .Z(\mreg/_06187_ ) );
BUF_X1 \mreg/_13177_ ( .A(\mreg/_00317_ ), .Z(\mreg/_06188_ ) );
BUF_X1 \mreg/_13178_ ( .A(\mreg/_00318_ ), .Z(\mreg/_06189_ ) );
BUF_X1 \mreg/_13179_ ( .A(\mreg/_00319_ ), .Z(\mreg/_06190_ ) );
BUF_X1 \mreg/_13180_ ( .A(\mreg/_00320_ ), .Z(\mreg/_06191_ ) );
BUF_X1 \mreg/_13181_ ( .A(\mreg/_00321_ ), .Z(\mreg/_06192_ ) );
BUF_X1 \mreg/_13182_ ( .A(\mreg/_00322_ ), .Z(\mreg/_06193_ ) );
BUF_X1 \mreg/_13183_ ( .A(\mreg/_00323_ ), .Z(\mreg/_06194_ ) );
BUF_X1 \mreg/_13184_ ( .A(\mreg/_00324_ ), .Z(\mreg/_06195_ ) );
BUF_X1 \mreg/_13185_ ( .A(\mreg/_00325_ ), .Z(\mreg/_06196_ ) );
BUF_X1 \mreg/_13186_ ( .A(\mreg/_00326_ ), .Z(\mreg/_06197_ ) );
BUF_X1 \mreg/_13187_ ( .A(\mreg/_00327_ ), .Z(\mreg/_06198_ ) );
BUF_X1 \mreg/_13188_ ( .A(\mreg/_00328_ ), .Z(\mreg/_06199_ ) );
BUF_X1 \mreg/_13189_ ( .A(\mreg/_00329_ ), .Z(\mreg/_06200_ ) );
BUF_X1 \mreg/_13190_ ( .A(\mreg/_00330_ ), .Z(\mreg/_06201_ ) );
BUF_X1 \mreg/_13191_ ( .A(\mreg/_00331_ ), .Z(\mreg/_06202_ ) );
BUF_X1 \mreg/_13192_ ( .A(\mreg/_00332_ ), .Z(\mreg/_06203_ ) );
BUF_X1 \mreg/_13193_ ( .A(\mreg/_00333_ ), .Z(\mreg/_06204_ ) );
BUF_X1 \mreg/_13194_ ( .A(\mreg/_00334_ ), .Z(\mreg/_06205_ ) );
BUF_X1 \mreg/_13195_ ( .A(\mreg/_00335_ ), .Z(\mreg/_06206_ ) );
BUF_X1 \mreg/_13196_ ( .A(\mreg/_00336_ ), .Z(\mreg/_06207_ ) );
BUF_X1 \mreg/_13197_ ( .A(\mreg/_00337_ ), .Z(\mreg/_06208_ ) );
BUF_X1 \mreg/_13198_ ( .A(\mreg/_00338_ ), .Z(\mreg/_06209_ ) );
BUF_X1 \mreg/_13199_ ( .A(\mreg/_00339_ ), .Z(\mreg/_06210_ ) );
BUF_X1 \mreg/_13200_ ( .A(\mreg/_00340_ ), .Z(\mreg/_06211_ ) );
BUF_X1 \mreg/_13201_ ( .A(\mreg/_00341_ ), .Z(\mreg/_06212_ ) );
BUF_X1 \mreg/_13202_ ( .A(\mreg/_00342_ ), .Z(\mreg/_06213_ ) );
BUF_X1 \mreg/_13203_ ( .A(\mreg/_00343_ ), .Z(\mreg/_06214_ ) );
BUF_X1 \mreg/_13204_ ( .A(\mreg/_00344_ ), .Z(\mreg/_06215_ ) );
BUF_X1 \mreg/_13205_ ( .A(\mreg/_00345_ ), .Z(\mreg/_06216_ ) );
BUF_X1 \mreg/_13206_ ( .A(\mreg/_00346_ ), .Z(\mreg/_06217_ ) );
BUF_X1 \mreg/_13207_ ( .A(\mreg/_00347_ ), .Z(\mreg/_06218_ ) );
BUF_X1 \mreg/_13208_ ( .A(\mreg/_00348_ ), .Z(\mreg/_06219_ ) );
BUF_X1 \mreg/_13209_ ( .A(\mreg/_00349_ ), .Z(\mreg/_06220_ ) );
BUF_X1 \mreg/_13210_ ( .A(\mreg/_00350_ ), .Z(\mreg/_06221_ ) );
BUF_X1 \mreg/_13211_ ( .A(\mreg/_00351_ ), .Z(\mreg/_06222_ ) );
BUF_X1 \mreg/_13212_ ( .A(\mreg/_00352_ ), .Z(\mreg/_06223_ ) );
BUF_X1 \mreg/_13213_ ( .A(\mreg/_00353_ ), .Z(\mreg/_06224_ ) );
BUF_X1 \mreg/_13214_ ( .A(\mreg/_00354_ ), .Z(\mreg/_06225_ ) );
BUF_X1 \mreg/_13215_ ( .A(\mreg/_00355_ ), .Z(\mreg/_06226_ ) );
BUF_X1 \mreg/_13216_ ( .A(\mreg/_00356_ ), .Z(\mreg/_06227_ ) );
BUF_X1 \mreg/_13217_ ( .A(\mreg/_00357_ ), .Z(\mreg/_06228_ ) );
BUF_X1 \mreg/_13218_ ( .A(\mreg/_00358_ ), .Z(\mreg/_06229_ ) );
BUF_X1 \mreg/_13219_ ( .A(\mreg/_00359_ ), .Z(\mreg/_06230_ ) );
BUF_X1 \mreg/_13220_ ( .A(\mreg/_00360_ ), .Z(\mreg/_06231_ ) );
BUF_X1 \mreg/_13221_ ( .A(\mreg/_00361_ ), .Z(\mreg/_06232_ ) );
BUF_X1 \mreg/_13222_ ( .A(\mreg/_00362_ ), .Z(\mreg/_06233_ ) );
BUF_X1 \mreg/_13223_ ( .A(\mreg/_00363_ ), .Z(\mreg/_06234_ ) );
BUF_X1 \mreg/_13224_ ( .A(\mreg/_00364_ ), .Z(\mreg/_06235_ ) );
BUF_X1 \mreg/_13225_ ( .A(\mreg/_00365_ ), .Z(\mreg/_06236_ ) );
BUF_X1 \mreg/_13226_ ( .A(\mreg/_00366_ ), .Z(\mreg/_06237_ ) );
BUF_X1 \mreg/_13227_ ( .A(\mreg/_00367_ ), .Z(\mreg/_06238_ ) );
BUF_X1 \mreg/_13228_ ( .A(\mreg/_00368_ ), .Z(\mreg/_06239_ ) );
BUF_X1 \mreg/_13229_ ( .A(\mreg/_00369_ ), .Z(\mreg/_06240_ ) );
BUF_X1 \mreg/_13230_ ( .A(\mreg/_00370_ ), .Z(\mreg/_06241_ ) );
BUF_X1 \mreg/_13231_ ( .A(\mreg/_00371_ ), .Z(\mreg/_06242_ ) );
BUF_X1 \mreg/_13232_ ( .A(\mreg/_00372_ ), .Z(\mreg/_06243_ ) );
BUF_X1 \mreg/_13233_ ( .A(\mreg/_00373_ ), .Z(\mreg/_06244_ ) );
BUF_X1 \mreg/_13234_ ( .A(\mreg/_00374_ ), .Z(\mreg/_06245_ ) );
BUF_X1 \mreg/_13235_ ( .A(\mreg/_00375_ ), .Z(\mreg/_06246_ ) );
BUF_X1 \mreg/_13236_ ( .A(\mreg/_00376_ ), .Z(\mreg/_06247_ ) );
BUF_X1 \mreg/_13237_ ( .A(\mreg/_00377_ ), .Z(\mreg/_06248_ ) );
BUF_X1 \mreg/_13238_ ( .A(\mreg/_00378_ ), .Z(\mreg/_06249_ ) );
BUF_X1 \mreg/_13239_ ( .A(\mreg/_00379_ ), .Z(\mreg/_06250_ ) );
BUF_X1 \mreg/_13240_ ( .A(\mreg/_00380_ ), .Z(\mreg/_06251_ ) );
BUF_X1 \mreg/_13241_ ( .A(\mreg/_00381_ ), .Z(\mreg/_06252_ ) );
BUF_X1 \mreg/_13242_ ( .A(\mreg/_00382_ ), .Z(\mreg/_06253_ ) );
BUF_X1 \mreg/_13243_ ( .A(\mreg/_00383_ ), .Z(\mreg/_06254_ ) );
BUF_X1 \mreg/_13244_ ( .A(\mreg/_00384_ ), .Z(\mreg/_06255_ ) );
BUF_X1 \mreg/_13245_ ( .A(\mreg/_00385_ ), .Z(\mreg/_06256_ ) );
BUF_X1 \mreg/_13246_ ( .A(\mreg/_00386_ ), .Z(\mreg/_06257_ ) );
BUF_X1 \mreg/_13247_ ( .A(\mreg/_00387_ ), .Z(\mreg/_06258_ ) );
BUF_X1 \mreg/_13248_ ( .A(\mreg/_00388_ ), .Z(\mreg/_06259_ ) );
BUF_X1 \mreg/_13249_ ( .A(\mreg/_00389_ ), .Z(\mreg/_06260_ ) );
BUF_X1 \mreg/_13250_ ( .A(\mreg/_00390_ ), .Z(\mreg/_06261_ ) );
BUF_X1 \mreg/_13251_ ( .A(\mreg/_00391_ ), .Z(\mreg/_06262_ ) );
BUF_X1 \mreg/_13252_ ( .A(\mreg/_00392_ ), .Z(\mreg/_06263_ ) );
BUF_X1 \mreg/_13253_ ( .A(\mreg/_00393_ ), .Z(\mreg/_06264_ ) );
BUF_X1 \mreg/_13254_ ( .A(\mreg/_00394_ ), .Z(\mreg/_06265_ ) );
BUF_X1 \mreg/_13255_ ( .A(\mreg/_00395_ ), .Z(\mreg/_06266_ ) );
BUF_X1 \mreg/_13256_ ( .A(\mreg/_00396_ ), .Z(\mreg/_06267_ ) );
BUF_X1 \mreg/_13257_ ( .A(\mreg/_00397_ ), .Z(\mreg/_06268_ ) );
BUF_X1 \mreg/_13258_ ( .A(\mreg/_00398_ ), .Z(\mreg/_06269_ ) );
BUF_X1 \mreg/_13259_ ( .A(\mreg/_00399_ ), .Z(\mreg/_06270_ ) );
BUF_X1 \mreg/_13260_ ( .A(\mreg/_00400_ ), .Z(\mreg/_06271_ ) );
BUF_X1 \mreg/_13261_ ( .A(\mreg/_00401_ ), .Z(\mreg/_06272_ ) );
BUF_X1 \mreg/_13262_ ( .A(\mreg/_00402_ ), .Z(\mreg/_06273_ ) );
BUF_X1 \mreg/_13263_ ( .A(\mreg/_00403_ ), .Z(\mreg/_06274_ ) );
BUF_X1 \mreg/_13264_ ( .A(\mreg/_00404_ ), .Z(\mreg/_06275_ ) );
BUF_X1 \mreg/_13265_ ( .A(\mreg/_00405_ ), .Z(\mreg/_06276_ ) );
BUF_X1 \mreg/_13266_ ( .A(\mreg/_00406_ ), .Z(\mreg/_06277_ ) );
BUF_X1 \mreg/_13267_ ( .A(\mreg/_00407_ ), .Z(\mreg/_06278_ ) );
BUF_X1 \mreg/_13268_ ( .A(\mreg/_00408_ ), .Z(\mreg/_06279_ ) );
BUF_X1 \mreg/_13269_ ( .A(\mreg/_00409_ ), .Z(\mreg/_06280_ ) );
BUF_X1 \mreg/_13270_ ( .A(\mreg/_00410_ ), .Z(\mreg/_06281_ ) );
BUF_X1 \mreg/_13271_ ( .A(\mreg/_00411_ ), .Z(\mreg/_06282_ ) );
BUF_X1 \mreg/_13272_ ( .A(\mreg/_00412_ ), .Z(\mreg/_06283_ ) );
BUF_X1 \mreg/_13273_ ( .A(\mreg/_00413_ ), .Z(\mreg/_06284_ ) );
BUF_X1 \mreg/_13274_ ( .A(\mreg/_00414_ ), .Z(\mreg/_06285_ ) );
BUF_X1 \mreg/_13275_ ( .A(\mreg/_00415_ ), .Z(\mreg/_06286_ ) );
BUF_X1 \mreg/_13276_ ( .A(\mreg/_00416_ ), .Z(\mreg/_06287_ ) );
BUF_X1 \mreg/_13277_ ( .A(\mreg/_00417_ ), .Z(\mreg/_06288_ ) );
BUF_X1 \mreg/_13278_ ( .A(\mreg/_00418_ ), .Z(\mreg/_06289_ ) );
BUF_X1 \mreg/_13279_ ( .A(\mreg/_00419_ ), .Z(\mreg/_06290_ ) );
BUF_X1 \mreg/_13280_ ( .A(\mreg/_00420_ ), .Z(\mreg/_06291_ ) );
BUF_X1 \mreg/_13281_ ( .A(\mreg/_00421_ ), .Z(\mreg/_06292_ ) );
BUF_X1 \mreg/_13282_ ( .A(\mreg/_00422_ ), .Z(\mreg/_06293_ ) );
BUF_X1 \mreg/_13283_ ( .A(\mreg/_00423_ ), .Z(\mreg/_06294_ ) );
BUF_X1 \mreg/_13284_ ( .A(\mreg/_00424_ ), .Z(\mreg/_06295_ ) );
BUF_X1 \mreg/_13285_ ( .A(\mreg/_00425_ ), .Z(\mreg/_06296_ ) );
BUF_X1 \mreg/_13286_ ( .A(\mreg/_00426_ ), .Z(\mreg/_06297_ ) );
BUF_X1 \mreg/_13287_ ( .A(\mreg/_00427_ ), .Z(\mreg/_06298_ ) );
BUF_X1 \mreg/_13288_ ( .A(\mreg/_00428_ ), .Z(\mreg/_06299_ ) );
BUF_X1 \mreg/_13289_ ( .A(\mreg/_00429_ ), .Z(\mreg/_06300_ ) );
BUF_X1 \mreg/_13290_ ( .A(\mreg/_00430_ ), .Z(\mreg/_06301_ ) );
BUF_X1 \mreg/_13291_ ( .A(\mreg/_00431_ ), .Z(\mreg/_06302_ ) );
BUF_X1 \mreg/_13292_ ( .A(\mreg/_00432_ ), .Z(\mreg/_06303_ ) );
BUF_X1 \mreg/_13293_ ( .A(\mreg/_00433_ ), .Z(\mreg/_06304_ ) );
BUF_X1 \mreg/_13294_ ( .A(\mreg/_00434_ ), .Z(\mreg/_06305_ ) );
BUF_X1 \mreg/_13295_ ( .A(\mreg/_00435_ ), .Z(\mreg/_06306_ ) );
BUF_X1 \mreg/_13296_ ( .A(\mreg/_00436_ ), .Z(\mreg/_06307_ ) );
BUF_X1 \mreg/_13297_ ( .A(\mreg/_00437_ ), .Z(\mreg/_06308_ ) );
BUF_X1 \mreg/_13298_ ( .A(\mreg/_00438_ ), .Z(\mreg/_06309_ ) );
BUF_X1 \mreg/_13299_ ( .A(\mreg/_00439_ ), .Z(\mreg/_06310_ ) );
BUF_X1 \mreg/_13300_ ( .A(\mreg/_00440_ ), .Z(\mreg/_06311_ ) );
BUF_X1 \mreg/_13301_ ( .A(\mreg/_00441_ ), .Z(\mreg/_06312_ ) );
BUF_X1 \mreg/_13302_ ( .A(\mreg/_00442_ ), .Z(\mreg/_06313_ ) );
BUF_X1 \mreg/_13303_ ( .A(\mreg/_00443_ ), .Z(\mreg/_06314_ ) );
BUF_X1 \mreg/_13304_ ( .A(\mreg/_00444_ ), .Z(\mreg/_06315_ ) );
BUF_X1 \mreg/_13305_ ( .A(\mreg/_00445_ ), .Z(\mreg/_06316_ ) );
BUF_X1 \mreg/_13306_ ( .A(\mreg/_00446_ ), .Z(\mreg/_06317_ ) );
BUF_X1 \mreg/_13307_ ( .A(\mreg/_00447_ ), .Z(\mreg/_06318_ ) );
BUF_X1 \mreg/_13308_ ( .A(\mreg/_00448_ ), .Z(\mreg/_06319_ ) );
BUF_X1 \mreg/_13309_ ( .A(\mreg/_00449_ ), .Z(\mreg/_06320_ ) );
BUF_X1 \mreg/_13310_ ( .A(\mreg/_00450_ ), .Z(\mreg/_06321_ ) );
BUF_X1 \mreg/_13311_ ( .A(\mreg/_00451_ ), .Z(\mreg/_06322_ ) );
BUF_X1 \mreg/_13312_ ( .A(\mreg/_00452_ ), .Z(\mreg/_06323_ ) );
BUF_X1 \mreg/_13313_ ( .A(\mreg/_00453_ ), .Z(\mreg/_06324_ ) );
BUF_X1 \mreg/_13314_ ( .A(\mreg/_00454_ ), .Z(\mreg/_06325_ ) );
BUF_X1 \mreg/_13315_ ( .A(\mreg/_00455_ ), .Z(\mreg/_06326_ ) );
BUF_X1 \mreg/_13316_ ( .A(\mreg/_00456_ ), .Z(\mreg/_06327_ ) );
BUF_X1 \mreg/_13317_ ( .A(\mreg/_00457_ ), .Z(\mreg/_06328_ ) );
BUF_X1 \mreg/_13318_ ( .A(\mreg/_00458_ ), .Z(\mreg/_06329_ ) );
BUF_X1 \mreg/_13319_ ( .A(\mreg/_00459_ ), .Z(\mreg/_06330_ ) );
BUF_X1 \mreg/_13320_ ( .A(\mreg/_00460_ ), .Z(\mreg/_06331_ ) );
BUF_X1 \mreg/_13321_ ( .A(\mreg/_00461_ ), .Z(\mreg/_06332_ ) );
BUF_X1 \mreg/_13322_ ( .A(\mreg/_00462_ ), .Z(\mreg/_06333_ ) );
BUF_X1 \mreg/_13323_ ( .A(\mreg/_00463_ ), .Z(\mreg/_06334_ ) );
BUF_X1 \mreg/_13324_ ( .A(\mreg/_00464_ ), .Z(\mreg/_06335_ ) );
BUF_X1 \mreg/_13325_ ( .A(\mreg/_00465_ ), .Z(\mreg/_06336_ ) );
BUF_X1 \mreg/_13326_ ( .A(\mreg/_00466_ ), .Z(\mreg/_06337_ ) );
BUF_X1 \mreg/_13327_ ( .A(\mreg/_00467_ ), .Z(\mreg/_06338_ ) );
BUF_X1 \mreg/_13328_ ( .A(\mreg/_00468_ ), .Z(\mreg/_06339_ ) );
BUF_X1 \mreg/_13329_ ( .A(\mreg/_00469_ ), .Z(\mreg/_06340_ ) );
BUF_X1 \mreg/_13330_ ( .A(\mreg/_00470_ ), .Z(\mreg/_06341_ ) );
BUF_X1 \mreg/_13331_ ( .A(\mreg/_00471_ ), .Z(\mreg/_06342_ ) );
BUF_X1 \mreg/_13332_ ( .A(\mreg/_00472_ ), .Z(\mreg/_06343_ ) );
BUF_X1 \mreg/_13333_ ( .A(\mreg/_00473_ ), .Z(\mreg/_06344_ ) );
BUF_X1 \mreg/_13334_ ( .A(\mreg/_00474_ ), .Z(\mreg/_06345_ ) );
BUF_X1 \mreg/_13335_ ( .A(\mreg/_00475_ ), .Z(\mreg/_06346_ ) );
BUF_X1 \mreg/_13336_ ( .A(\mreg/_00476_ ), .Z(\mreg/_06347_ ) );
BUF_X1 \mreg/_13337_ ( .A(\mreg/_00477_ ), .Z(\mreg/_06348_ ) );
BUF_X1 \mreg/_13338_ ( .A(\mreg/_00478_ ), .Z(\mreg/_06349_ ) );
BUF_X1 \mreg/_13339_ ( .A(\mreg/_00479_ ), .Z(\mreg/_06350_ ) );
BUF_X1 \mreg/_13340_ ( .A(\mreg/_00480_ ), .Z(\mreg/_06351_ ) );
BUF_X1 \mreg/_13341_ ( .A(\mreg/_00481_ ), .Z(\mreg/_06352_ ) );
BUF_X1 \mreg/_13342_ ( .A(\mreg/_00482_ ), .Z(\mreg/_06353_ ) );
BUF_X1 \mreg/_13343_ ( .A(\mreg/_00483_ ), .Z(\mreg/_06354_ ) );
BUF_X1 \mreg/_13344_ ( .A(\mreg/_00484_ ), .Z(\mreg/_06355_ ) );
BUF_X1 \mreg/_13345_ ( .A(\mreg/_00485_ ), .Z(\mreg/_06356_ ) );
BUF_X1 \mreg/_13346_ ( .A(\mreg/_00486_ ), .Z(\mreg/_06357_ ) );
BUF_X1 \mreg/_13347_ ( .A(\mreg/_00487_ ), .Z(\mreg/_06358_ ) );
BUF_X1 \mreg/_13348_ ( .A(\mreg/_00488_ ), .Z(\mreg/_06359_ ) );
BUF_X1 \mreg/_13349_ ( .A(\mreg/_00489_ ), .Z(\mreg/_06360_ ) );
BUF_X1 \mreg/_13350_ ( .A(\mreg/_00490_ ), .Z(\mreg/_06361_ ) );
BUF_X1 \mreg/_13351_ ( .A(\mreg/_00491_ ), .Z(\mreg/_06362_ ) );
BUF_X1 \mreg/_13352_ ( .A(\mreg/_00492_ ), .Z(\mreg/_06363_ ) );
BUF_X1 \mreg/_13353_ ( .A(\mreg/_00493_ ), .Z(\mreg/_06364_ ) );
BUF_X1 \mreg/_13354_ ( .A(\mreg/_00494_ ), .Z(\mreg/_06365_ ) );
BUF_X1 \mreg/_13355_ ( .A(\mreg/_00495_ ), .Z(\mreg/_06366_ ) );
BUF_X1 \mreg/_13356_ ( .A(\mreg/_00496_ ), .Z(\mreg/_06367_ ) );
BUF_X1 \mreg/_13357_ ( .A(\mreg/_00497_ ), .Z(\mreg/_06368_ ) );
BUF_X1 \mreg/_13358_ ( .A(\mreg/_00498_ ), .Z(\mreg/_06369_ ) );
BUF_X1 \mreg/_13359_ ( .A(\mreg/_00499_ ), .Z(\mreg/_06370_ ) );
BUF_X1 \mreg/_13360_ ( .A(\mreg/_00500_ ), .Z(\mreg/_06371_ ) );
BUF_X1 \mreg/_13361_ ( .A(\mreg/_00501_ ), .Z(\mreg/_06372_ ) );
BUF_X1 \mreg/_13362_ ( .A(\mreg/_00502_ ), .Z(\mreg/_06373_ ) );
BUF_X1 \mreg/_13363_ ( .A(\mreg/_00503_ ), .Z(\mreg/_06374_ ) );
BUF_X1 \mreg/_13364_ ( .A(\mreg/_00504_ ), .Z(\mreg/_06375_ ) );
BUF_X1 \mreg/_13365_ ( .A(\mreg/_00505_ ), .Z(\mreg/_06376_ ) );
BUF_X1 \mreg/_13366_ ( .A(\mreg/_00506_ ), .Z(\mreg/_06377_ ) );
BUF_X1 \mreg/_13367_ ( .A(\mreg/_00507_ ), .Z(\mreg/_06378_ ) );
BUF_X1 \mreg/_13368_ ( .A(\mreg/_00508_ ), .Z(\mreg/_06379_ ) );
BUF_X1 \mreg/_13369_ ( .A(\mreg/_00509_ ), .Z(\mreg/_06380_ ) );
BUF_X1 \mreg/_13370_ ( .A(\mreg/_00510_ ), .Z(\mreg/_06381_ ) );
BUF_X1 \mreg/_13371_ ( .A(\mreg/_00511_ ), .Z(\mreg/_06382_ ) );
BUF_X1 \mreg/_13372_ ( .A(\mreg/_00512_ ), .Z(\mreg/_06383_ ) );
BUF_X1 \mreg/_13373_ ( .A(\mreg/_00513_ ), .Z(\mreg/_06384_ ) );
BUF_X1 \mreg/_13374_ ( .A(\mreg/_00514_ ), .Z(\mreg/_06385_ ) );
BUF_X1 \mreg/_13375_ ( .A(\mreg/_00515_ ), .Z(\mreg/_06386_ ) );
BUF_X1 \mreg/_13376_ ( .A(\mreg/_00516_ ), .Z(\mreg/_06387_ ) );
BUF_X1 \mreg/_13377_ ( .A(\mreg/_00517_ ), .Z(\mreg/_06388_ ) );
BUF_X1 \mreg/_13378_ ( .A(\mreg/_00518_ ), .Z(\mreg/_06389_ ) );
BUF_X1 \mreg/_13379_ ( .A(\mreg/_00519_ ), .Z(\mreg/_06390_ ) );
BUF_X1 \mreg/_13380_ ( .A(\mreg/_00520_ ), .Z(\mreg/_06391_ ) );
BUF_X1 \mreg/_13381_ ( .A(\mreg/_00521_ ), .Z(\mreg/_06392_ ) );
BUF_X1 \mreg/_13382_ ( .A(\mreg/_00522_ ), .Z(\mreg/_06393_ ) );
BUF_X1 \mreg/_13383_ ( .A(\mreg/_00523_ ), .Z(\mreg/_06394_ ) );
BUF_X1 \mreg/_13384_ ( .A(\mreg/_00524_ ), .Z(\mreg/_06395_ ) );
BUF_X1 \mreg/_13385_ ( .A(\mreg/_00525_ ), .Z(\mreg/_06396_ ) );
BUF_X1 \mreg/_13386_ ( .A(\mreg/_00526_ ), .Z(\mreg/_06397_ ) );
BUF_X1 \mreg/_13387_ ( .A(\mreg/_00527_ ), .Z(\mreg/_06398_ ) );
BUF_X1 \mreg/_13388_ ( .A(\mreg/_00528_ ), .Z(\mreg/_06399_ ) );
BUF_X1 \mreg/_13389_ ( .A(\mreg/_00529_ ), .Z(\mreg/_06400_ ) );
BUF_X1 \mreg/_13390_ ( .A(\mreg/_00530_ ), .Z(\mreg/_06401_ ) );
BUF_X1 \mreg/_13391_ ( .A(\mreg/_00531_ ), .Z(\mreg/_06402_ ) );
BUF_X1 \mreg/_13392_ ( .A(\mreg/_00532_ ), .Z(\mreg/_06403_ ) );
BUF_X1 \mreg/_13393_ ( .A(\mreg/_00533_ ), .Z(\mreg/_06404_ ) );
BUF_X1 \mreg/_13394_ ( .A(\mreg/_00534_ ), .Z(\mreg/_06405_ ) );
BUF_X1 \mreg/_13395_ ( .A(\mreg/_00535_ ), .Z(\mreg/_06406_ ) );
BUF_X1 \mreg/_13396_ ( .A(\mreg/_00536_ ), .Z(\mreg/_06407_ ) );
BUF_X1 \mreg/_13397_ ( .A(\mreg/_00537_ ), .Z(\mreg/_06408_ ) );
BUF_X1 \mreg/_13398_ ( .A(\mreg/_00538_ ), .Z(\mreg/_06409_ ) );
BUF_X1 \mreg/_13399_ ( .A(\mreg/_00539_ ), .Z(\mreg/_06410_ ) );
BUF_X1 \mreg/_13400_ ( .A(\mreg/_00540_ ), .Z(\mreg/_06411_ ) );
BUF_X1 \mreg/_13401_ ( .A(\mreg/_00541_ ), .Z(\mreg/_06412_ ) );
BUF_X1 \mreg/_13402_ ( .A(\mreg/_00542_ ), .Z(\mreg/_06413_ ) );
BUF_X1 \mreg/_13403_ ( .A(\mreg/_00543_ ), .Z(\mreg/_06414_ ) );
BUF_X1 \mreg/_13404_ ( .A(\mreg/_00544_ ), .Z(\mreg/_06415_ ) );
BUF_X1 \mreg/_13405_ ( .A(\mreg/_00545_ ), .Z(\mreg/_06416_ ) );
BUF_X1 \mreg/_13406_ ( .A(\mreg/_00546_ ), .Z(\mreg/_06417_ ) );
BUF_X1 \mreg/_13407_ ( .A(\mreg/_00547_ ), .Z(\mreg/_06418_ ) );
BUF_X1 \mreg/_13408_ ( .A(\mreg/_00548_ ), .Z(\mreg/_06419_ ) );
BUF_X1 \mreg/_13409_ ( .A(\mreg/_00549_ ), .Z(\mreg/_06420_ ) );
BUF_X1 \mreg/_13410_ ( .A(\mreg/_00550_ ), .Z(\mreg/_06421_ ) );
BUF_X1 \mreg/_13411_ ( .A(\mreg/_00551_ ), .Z(\mreg/_06422_ ) );
BUF_X1 \mreg/_13412_ ( .A(\mreg/_00552_ ), .Z(\mreg/_06423_ ) );
BUF_X1 \mreg/_13413_ ( .A(\mreg/_00553_ ), .Z(\mreg/_06424_ ) );
BUF_X1 \mreg/_13414_ ( .A(\mreg/_00554_ ), .Z(\mreg/_06425_ ) );
BUF_X1 \mreg/_13415_ ( .A(\mreg/_00555_ ), .Z(\mreg/_06426_ ) );
BUF_X1 \mreg/_13416_ ( .A(\mreg/_00556_ ), .Z(\mreg/_06427_ ) );
BUF_X1 \mreg/_13417_ ( .A(\mreg/_00557_ ), .Z(\mreg/_06428_ ) );
BUF_X1 \mreg/_13418_ ( .A(\mreg/_00558_ ), .Z(\mreg/_06429_ ) );
BUF_X1 \mreg/_13419_ ( .A(\mreg/_00559_ ), .Z(\mreg/_06430_ ) );
BUF_X1 \mreg/_13420_ ( .A(\mreg/_00560_ ), .Z(\mreg/_06431_ ) );
BUF_X1 \mreg/_13421_ ( .A(\mreg/_00561_ ), .Z(\mreg/_06432_ ) );
BUF_X1 \mreg/_13422_ ( .A(\mreg/_00562_ ), .Z(\mreg/_06433_ ) );
BUF_X1 \mreg/_13423_ ( .A(\mreg/_00563_ ), .Z(\mreg/_06434_ ) );
BUF_X1 \mreg/_13424_ ( .A(\mreg/_00564_ ), .Z(\mreg/_06435_ ) );
BUF_X1 \mreg/_13425_ ( .A(\mreg/_00565_ ), .Z(\mreg/_06436_ ) );
BUF_X1 \mreg/_13426_ ( .A(\mreg/_00566_ ), .Z(\mreg/_06437_ ) );
BUF_X1 \mreg/_13427_ ( .A(\mreg/_00567_ ), .Z(\mreg/_06438_ ) );
BUF_X1 \mreg/_13428_ ( .A(\mreg/_00568_ ), .Z(\mreg/_06439_ ) );
BUF_X1 \mreg/_13429_ ( .A(\mreg/_00569_ ), .Z(\mreg/_06440_ ) );
BUF_X1 \mreg/_13430_ ( .A(\mreg/_00570_ ), .Z(\mreg/_06441_ ) );
BUF_X1 \mreg/_13431_ ( .A(\mreg/_00571_ ), .Z(\mreg/_06442_ ) );
BUF_X1 \mreg/_13432_ ( .A(\mreg/_00572_ ), .Z(\mreg/_06443_ ) );
BUF_X1 \mreg/_13433_ ( .A(\mreg/_00573_ ), .Z(\mreg/_06444_ ) );
BUF_X1 \mreg/_13434_ ( .A(\mreg/_00574_ ), .Z(\mreg/_06445_ ) );
BUF_X1 \mreg/_13435_ ( .A(\mreg/_00575_ ), .Z(\mreg/_06446_ ) );
BUF_X1 \mreg/_13436_ ( .A(\mreg/_00576_ ), .Z(\mreg/_06447_ ) );
BUF_X1 \mreg/_13437_ ( .A(\mreg/_00577_ ), .Z(\mreg/_06448_ ) );
BUF_X1 \mreg/_13438_ ( .A(\mreg/_00578_ ), .Z(\mreg/_06449_ ) );
BUF_X1 \mreg/_13439_ ( .A(\mreg/_00579_ ), .Z(\mreg/_06450_ ) );
BUF_X1 \mreg/_13440_ ( .A(\mreg/_00580_ ), .Z(\mreg/_06451_ ) );
BUF_X1 \mreg/_13441_ ( .A(\mreg/_00581_ ), .Z(\mreg/_06452_ ) );
BUF_X1 \mreg/_13442_ ( .A(\mreg/_00582_ ), .Z(\mreg/_06453_ ) );
BUF_X1 \mreg/_13443_ ( .A(\mreg/_00583_ ), .Z(\mreg/_06454_ ) );
BUF_X1 \mreg/_13444_ ( .A(\mreg/_00584_ ), .Z(\mreg/_06455_ ) );
BUF_X1 \mreg/_13445_ ( .A(\mreg/_00585_ ), .Z(\mreg/_06456_ ) );
BUF_X1 \mreg/_13446_ ( .A(\mreg/_00586_ ), .Z(\mreg/_06457_ ) );
BUF_X1 \mreg/_13447_ ( .A(\mreg/_00587_ ), .Z(\mreg/_06458_ ) );
BUF_X1 \mreg/_13448_ ( .A(\mreg/_00588_ ), .Z(\mreg/_06459_ ) );
BUF_X1 \mreg/_13449_ ( .A(\mreg/_00589_ ), .Z(\mreg/_06460_ ) );
BUF_X1 \mreg/_13450_ ( .A(\mreg/_00590_ ), .Z(\mreg/_06461_ ) );
BUF_X1 \mreg/_13451_ ( .A(\mreg/_00591_ ), .Z(\mreg/_06462_ ) );
BUF_X1 \mreg/_13452_ ( .A(\mreg/_00592_ ), .Z(\mreg/_06463_ ) );
BUF_X1 \mreg/_13453_ ( .A(\mreg/_00593_ ), .Z(\mreg/_06464_ ) );
BUF_X1 \mreg/_13454_ ( .A(\mreg/_00594_ ), .Z(\mreg/_06465_ ) );
BUF_X1 \mreg/_13455_ ( .A(\mreg/_00595_ ), .Z(\mreg/_06466_ ) );
BUF_X1 \mreg/_13456_ ( .A(\mreg/_00596_ ), .Z(\mreg/_06467_ ) );
BUF_X1 \mreg/_13457_ ( .A(\mreg/_00597_ ), .Z(\mreg/_06468_ ) );
BUF_X1 \mreg/_13458_ ( .A(\mreg/_00598_ ), .Z(\mreg/_06469_ ) );
BUF_X1 \mreg/_13459_ ( .A(\mreg/_00599_ ), .Z(\mreg/_06470_ ) );
BUF_X1 \mreg/_13460_ ( .A(\mreg/_00600_ ), .Z(\mreg/_06471_ ) );
BUF_X1 \mreg/_13461_ ( .A(\mreg/_00601_ ), .Z(\mreg/_06472_ ) );
BUF_X1 \mreg/_13462_ ( .A(\mreg/_00602_ ), .Z(\mreg/_06473_ ) );
BUF_X1 \mreg/_13463_ ( .A(\mreg/_00603_ ), .Z(\mreg/_06474_ ) );
BUF_X1 \mreg/_13464_ ( .A(\mreg/_00604_ ), .Z(\mreg/_06475_ ) );
BUF_X1 \mreg/_13465_ ( .A(\mreg/_00605_ ), .Z(\mreg/_06476_ ) );
BUF_X1 \mreg/_13466_ ( .A(\mreg/_00606_ ), .Z(\mreg/_06477_ ) );
BUF_X1 \mreg/_13467_ ( .A(\mreg/_00607_ ), .Z(\mreg/_06478_ ) );
BUF_X1 \mreg/_13468_ ( .A(\mreg/_00608_ ), .Z(\mreg/_06479_ ) );
BUF_X1 \mreg/_13469_ ( .A(\mreg/_00609_ ), .Z(\mreg/_06480_ ) );
BUF_X1 \mreg/_13470_ ( .A(\mreg/_00610_ ), .Z(\mreg/_06481_ ) );
BUF_X1 \mreg/_13471_ ( .A(\mreg/_00611_ ), .Z(\mreg/_06482_ ) );
BUF_X1 \mreg/_13472_ ( .A(\mreg/_00612_ ), .Z(\mreg/_06483_ ) );
BUF_X1 \mreg/_13473_ ( .A(\mreg/_00613_ ), .Z(\mreg/_06484_ ) );
BUF_X1 \mreg/_13474_ ( .A(\mreg/_00614_ ), .Z(\mreg/_06485_ ) );
BUF_X1 \mreg/_13475_ ( .A(\mreg/_00615_ ), .Z(\mreg/_06486_ ) );
BUF_X1 \mreg/_13476_ ( .A(\mreg/_00616_ ), .Z(\mreg/_06487_ ) );
BUF_X1 \mreg/_13477_ ( .A(\mreg/_00617_ ), .Z(\mreg/_06488_ ) );
BUF_X1 \mreg/_13478_ ( .A(\mreg/_00618_ ), .Z(\mreg/_06489_ ) );
BUF_X1 \mreg/_13479_ ( .A(\mreg/_00619_ ), .Z(\mreg/_06490_ ) );
BUF_X1 \mreg/_13480_ ( .A(\mreg/_00620_ ), .Z(\mreg/_06491_ ) );
BUF_X1 \mreg/_13481_ ( .A(\mreg/_00621_ ), .Z(\mreg/_06492_ ) );
BUF_X1 \mreg/_13482_ ( .A(\mreg/_00622_ ), .Z(\mreg/_06493_ ) );
BUF_X1 \mreg/_13483_ ( .A(\mreg/_00623_ ), .Z(\mreg/_06494_ ) );
BUF_X1 \mreg/_13484_ ( .A(\mreg/_00624_ ), .Z(\mreg/_06495_ ) );
BUF_X1 \mreg/_13485_ ( .A(\mreg/_00625_ ), .Z(\mreg/_06496_ ) );
BUF_X1 \mreg/_13486_ ( .A(\mreg/_00626_ ), .Z(\mreg/_06497_ ) );
BUF_X1 \mreg/_13487_ ( .A(\mreg/_00627_ ), .Z(\mreg/_06498_ ) );
BUF_X1 \mreg/_13488_ ( .A(\mreg/_00628_ ), .Z(\mreg/_06499_ ) );
BUF_X1 \mreg/_13489_ ( .A(\mreg/_00629_ ), .Z(\mreg/_06500_ ) );
BUF_X1 \mreg/_13490_ ( .A(\mreg/_00630_ ), .Z(\mreg/_06501_ ) );
BUF_X1 \mreg/_13491_ ( .A(\mreg/_00631_ ), .Z(\mreg/_06502_ ) );
BUF_X1 \mreg/_13492_ ( .A(\mreg/_00632_ ), .Z(\mreg/_06503_ ) );
BUF_X1 \mreg/_13493_ ( .A(\mreg/_00633_ ), .Z(\mreg/_06504_ ) );
BUF_X1 \mreg/_13494_ ( .A(\mreg/_00634_ ), .Z(\mreg/_06505_ ) );
BUF_X1 \mreg/_13495_ ( .A(\mreg/_00635_ ), .Z(\mreg/_06506_ ) );
BUF_X1 \mreg/_13496_ ( .A(\mreg/_00636_ ), .Z(\mreg/_06507_ ) );
BUF_X1 \mreg/_13497_ ( .A(\mreg/_00637_ ), .Z(\mreg/_06508_ ) );
BUF_X1 \mreg/_13498_ ( .A(\mreg/_00638_ ), .Z(\mreg/_06509_ ) );
BUF_X1 \mreg/_13499_ ( .A(\mreg/_00639_ ), .Z(\mreg/_06510_ ) );
BUF_X1 \mreg/_13500_ ( .A(\mreg/_00640_ ), .Z(\mreg/_06511_ ) );
BUF_X1 \mreg/_13501_ ( .A(\mreg/_00641_ ), .Z(\mreg/_06512_ ) );
BUF_X1 \mreg/_13502_ ( .A(\mreg/_00642_ ), .Z(\mreg/_06513_ ) );
BUF_X1 \mreg/_13503_ ( .A(\mreg/_00643_ ), .Z(\mreg/_06514_ ) );
BUF_X1 \mreg/_13504_ ( .A(\mreg/_00644_ ), .Z(\mreg/_06515_ ) );
BUF_X1 \mreg/_13505_ ( .A(\mreg/_00645_ ), .Z(\mreg/_06516_ ) );
BUF_X1 \mreg/_13506_ ( .A(\mreg/_00646_ ), .Z(\mreg/_06517_ ) );
BUF_X1 \mreg/_13507_ ( .A(\mreg/_00647_ ), .Z(\mreg/_06518_ ) );
BUF_X1 \mreg/_13508_ ( .A(\mreg/_00648_ ), .Z(\mreg/_06519_ ) );
BUF_X1 \mreg/_13509_ ( .A(\mreg/_00649_ ), .Z(\mreg/_06520_ ) );
BUF_X1 \mreg/_13510_ ( .A(\mreg/_00650_ ), .Z(\mreg/_06521_ ) );
BUF_X1 \mreg/_13511_ ( .A(\mreg/_00651_ ), .Z(\mreg/_06522_ ) );
BUF_X1 \mreg/_13512_ ( .A(\mreg/_00652_ ), .Z(\mreg/_06523_ ) );
BUF_X1 \mreg/_13513_ ( .A(\mreg/_00653_ ), .Z(\mreg/_06524_ ) );
BUF_X1 \mreg/_13514_ ( .A(\mreg/_00654_ ), .Z(\mreg/_06525_ ) );
BUF_X1 \mreg/_13515_ ( .A(\mreg/_00655_ ), .Z(\mreg/_06526_ ) );
BUF_X1 \mreg/_13516_ ( .A(\mreg/_00656_ ), .Z(\mreg/_06527_ ) );
BUF_X1 \mreg/_13517_ ( .A(\mreg/_00657_ ), .Z(\mreg/_06528_ ) );
BUF_X1 \mreg/_13518_ ( .A(\mreg/_00658_ ), .Z(\mreg/_06529_ ) );
BUF_X1 \mreg/_13519_ ( .A(\mreg/_00659_ ), .Z(\mreg/_06530_ ) );
BUF_X1 \mreg/_13520_ ( .A(\mreg/_00660_ ), .Z(\mreg/_06531_ ) );
BUF_X1 \mreg/_13521_ ( .A(\mreg/_00661_ ), .Z(\mreg/_06532_ ) );
BUF_X1 \mreg/_13522_ ( .A(\mreg/_00662_ ), .Z(\mreg/_06533_ ) );
BUF_X1 \mreg/_13523_ ( .A(\mreg/_00663_ ), .Z(\mreg/_06534_ ) );
BUF_X1 \mreg/_13524_ ( .A(\mreg/_00664_ ), .Z(\mreg/_06535_ ) );
BUF_X1 \mreg/_13525_ ( .A(\mreg/_00665_ ), .Z(\mreg/_06536_ ) );
BUF_X1 \mreg/_13526_ ( .A(\mreg/_00666_ ), .Z(\mreg/_06537_ ) );
BUF_X1 \mreg/_13527_ ( .A(\mreg/_00667_ ), .Z(\mreg/_06538_ ) );
BUF_X1 \mreg/_13528_ ( .A(\mreg/_00668_ ), .Z(\mreg/_06539_ ) );
BUF_X1 \mreg/_13529_ ( .A(\mreg/_00669_ ), .Z(\mreg/_06540_ ) );
BUF_X1 \mreg/_13530_ ( .A(\mreg/_00670_ ), .Z(\mreg/_06541_ ) );
BUF_X1 \mreg/_13531_ ( .A(\mreg/_00671_ ), .Z(\mreg/_06542_ ) );
BUF_X1 \mreg/_13532_ ( .A(\mreg/_00672_ ), .Z(\mreg/_06543_ ) );
BUF_X1 \mreg/_13533_ ( .A(\mreg/_00673_ ), .Z(\mreg/_06544_ ) );
BUF_X1 \mreg/_13534_ ( .A(\mreg/_00674_ ), .Z(\mreg/_06545_ ) );
BUF_X1 \mreg/_13535_ ( .A(\mreg/_00675_ ), .Z(\mreg/_06546_ ) );
BUF_X1 \mreg/_13536_ ( .A(\mreg/_00676_ ), .Z(\mreg/_06547_ ) );
BUF_X1 \mreg/_13537_ ( .A(\mreg/_00677_ ), .Z(\mreg/_06548_ ) );
BUF_X1 \mreg/_13538_ ( .A(\mreg/_00678_ ), .Z(\mreg/_06549_ ) );
BUF_X1 \mreg/_13539_ ( .A(\mreg/_00679_ ), .Z(\mreg/_06550_ ) );
BUF_X1 \mreg/_13540_ ( .A(\mreg/_00680_ ), .Z(\mreg/_06551_ ) );
BUF_X1 \mreg/_13541_ ( .A(\mreg/_00681_ ), .Z(\mreg/_06552_ ) );
BUF_X1 \mreg/_13542_ ( .A(\mreg/_00682_ ), .Z(\mreg/_06553_ ) );
BUF_X1 \mreg/_13543_ ( .A(\mreg/_00683_ ), .Z(\mreg/_06554_ ) );
BUF_X1 \mreg/_13544_ ( .A(\mreg/_00684_ ), .Z(\mreg/_06555_ ) );
BUF_X1 \mreg/_13545_ ( .A(\mreg/_00685_ ), .Z(\mreg/_06556_ ) );
BUF_X1 \mreg/_13546_ ( .A(\mreg/_00686_ ), .Z(\mreg/_06557_ ) );
BUF_X1 \mreg/_13547_ ( .A(\mreg/_00687_ ), .Z(\mreg/_06558_ ) );
BUF_X1 \mreg/_13548_ ( .A(\mreg/_00688_ ), .Z(\mreg/_06559_ ) );
BUF_X1 \mreg/_13549_ ( .A(\mreg/_00689_ ), .Z(\mreg/_06560_ ) );
BUF_X1 \mreg/_13550_ ( .A(\mreg/_00690_ ), .Z(\mreg/_06561_ ) );
BUF_X1 \mreg/_13551_ ( .A(\mreg/_00691_ ), .Z(\mreg/_06562_ ) );
BUF_X1 \mreg/_13552_ ( .A(\mreg/_00692_ ), .Z(\mreg/_06563_ ) );
BUF_X1 \mreg/_13553_ ( .A(\mreg/_00693_ ), .Z(\mreg/_06564_ ) );
BUF_X1 \mreg/_13554_ ( .A(\mreg/_00694_ ), .Z(\mreg/_06565_ ) );
BUF_X1 \mreg/_13555_ ( .A(\mreg/_00695_ ), .Z(\mreg/_06566_ ) );
BUF_X1 \mreg/_13556_ ( .A(\mreg/_00696_ ), .Z(\mreg/_06567_ ) );
BUF_X1 \mreg/_13557_ ( .A(\mreg/_00697_ ), .Z(\mreg/_06568_ ) );
BUF_X1 \mreg/_13558_ ( .A(\mreg/_00698_ ), .Z(\mreg/_06569_ ) );
BUF_X1 \mreg/_13559_ ( .A(\mreg/_00699_ ), .Z(\mreg/_06570_ ) );
BUF_X1 \mreg/_13560_ ( .A(\mreg/_00700_ ), .Z(\mreg/_06571_ ) );
BUF_X1 \mreg/_13561_ ( .A(\mreg/_00701_ ), .Z(\mreg/_06572_ ) );
BUF_X1 \mreg/_13562_ ( .A(\mreg/_00702_ ), .Z(\mreg/_06573_ ) );
BUF_X1 \mreg/_13563_ ( .A(\mreg/_00703_ ), .Z(\mreg/_06574_ ) );
BUF_X1 \mreg/_13564_ ( .A(\mreg/_00704_ ), .Z(\mreg/_06575_ ) );
BUF_X1 \mreg/_13565_ ( .A(\mreg/_00705_ ), .Z(\mreg/_06576_ ) );
BUF_X1 \mreg/_13566_ ( .A(\mreg/_00706_ ), .Z(\mreg/_06577_ ) );
BUF_X1 \mreg/_13567_ ( .A(\mreg/_00707_ ), .Z(\mreg/_06578_ ) );
BUF_X1 \mreg/_13568_ ( .A(\mreg/_00708_ ), .Z(\mreg/_06579_ ) );
BUF_X1 \mreg/_13569_ ( .A(\mreg/_00709_ ), .Z(\mreg/_06580_ ) );
BUF_X1 \mreg/_13570_ ( .A(\mreg/_00710_ ), .Z(\mreg/_06581_ ) );
BUF_X1 \mreg/_13571_ ( .A(\mreg/_00711_ ), .Z(\mreg/_06582_ ) );
BUF_X1 \mreg/_13572_ ( .A(\mreg/_00712_ ), .Z(\mreg/_06583_ ) );
BUF_X1 \mreg/_13573_ ( .A(\mreg/_00713_ ), .Z(\mreg/_06584_ ) );
BUF_X1 \mreg/_13574_ ( .A(\mreg/_00714_ ), .Z(\mreg/_06585_ ) );
BUF_X1 \mreg/_13575_ ( .A(\mreg/_00715_ ), .Z(\mreg/_06586_ ) );
BUF_X1 \mreg/_13576_ ( .A(\mreg/_00716_ ), .Z(\mreg/_06587_ ) );
BUF_X1 \mreg/_13577_ ( .A(\mreg/_00717_ ), .Z(\mreg/_06588_ ) );
BUF_X1 \mreg/_13578_ ( .A(\mreg/_00718_ ), .Z(\mreg/_06589_ ) );
BUF_X1 \mreg/_13579_ ( .A(\mreg/_00719_ ), .Z(\mreg/_06590_ ) );
BUF_X1 \mreg/_13580_ ( .A(\mreg/_00720_ ), .Z(\mreg/_06591_ ) );
BUF_X1 \mreg/_13581_ ( .A(\mreg/_00721_ ), .Z(\mreg/_06592_ ) );
BUF_X1 \mreg/_13582_ ( .A(\mreg/_00722_ ), .Z(\mreg/_06593_ ) );
BUF_X1 \mreg/_13583_ ( .A(\mreg/_00723_ ), .Z(\mreg/_06594_ ) );
BUF_X1 \mreg/_13584_ ( .A(\mreg/_00724_ ), .Z(\mreg/_06595_ ) );
BUF_X1 \mreg/_13585_ ( .A(\mreg/_00725_ ), .Z(\mreg/_06596_ ) );
BUF_X1 \mreg/_13586_ ( .A(\mreg/_00726_ ), .Z(\mreg/_06597_ ) );
BUF_X1 \mreg/_13587_ ( .A(\mreg/_00727_ ), .Z(\mreg/_06598_ ) );
BUF_X1 \mreg/_13588_ ( .A(\mreg/_00728_ ), .Z(\mreg/_06599_ ) );
BUF_X1 \mreg/_13589_ ( .A(\mreg/_00729_ ), .Z(\mreg/_06600_ ) );
BUF_X1 \mreg/_13590_ ( .A(\mreg/_00730_ ), .Z(\mreg/_06601_ ) );
BUF_X1 \mreg/_13591_ ( .A(\mreg/_00731_ ), .Z(\mreg/_06602_ ) );
BUF_X1 \mreg/_13592_ ( .A(\mreg/_00732_ ), .Z(\mreg/_06603_ ) );
BUF_X1 \mreg/_13593_ ( .A(\mreg/_00733_ ), .Z(\mreg/_06604_ ) );
BUF_X1 \mreg/_13594_ ( .A(\mreg/_00734_ ), .Z(\mreg/_06605_ ) );
BUF_X1 \mreg/_13595_ ( .A(\mreg/_00735_ ), .Z(\mreg/_06606_ ) );
BUF_X1 \mreg/_13596_ ( .A(\mreg/_00736_ ), .Z(\mreg/_06607_ ) );
BUF_X1 \mreg/_13597_ ( .A(\mreg/_00737_ ), .Z(\mreg/_06608_ ) );
BUF_X1 \mreg/_13598_ ( .A(\mreg/_00738_ ), .Z(\mreg/_06609_ ) );
BUF_X1 \mreg/_13599_ ( .A(\mreg/_00739_ ), .Z(\mreg/_06610_ ) );
BUF_X1 \mreg/_13600_ ( .A(\mreg/_00740_ ), .Z(\mreg/_06611_ ) );
BUF_X1 \mreg/_13601_ ( .A(\mreg/_00741_ ), .Z(\mreg/_06612_ ) );
BUF_X1 \mreg/_13602_ ( .A(\mreg/_00742_ ), .Z(\mreg/_06613_ ) );
BUF_X1 \mreg/_13603_ ( .A(\mreg/_00743_ ), .Z(\mreg/_06614_ ) );
BUF_X1 \mreg/_13604_ ( .A(\mreg/_00744_ ), .Z(\mreg/_06615_ ) );
BUF_X1 \mreg/_13605_ ( .A(\mreg/_00745_ ), .Z(\mreg/_06616_ ) );
BUF_X1 \mreg/_13606_ ( .A(\mreg/_00746_ ), .Z(\mreg/_06617_ ) );
BUF_X1 \mreg/_13607_ ( .A(\mreg/_00747_ ), .Z(\mreg/_06618_ ) );
BUF_X1 \mreg/_13608_ ( .A(\mreg/_00748_ ), .Z(\mreg/_06619_ ) );
BUF_X1 \mreg/_13609_ ( .A(\mreg/_00749_ ), .Z(\mreg/_06620_ ) );
BUF_X1 \mreg/_13610_ ( .A(\mreg/_00750_ ), .Z(\mreg/_06621_ ) );
BUF_X1 \mreg/_13611_ ( .A(\mreg/_00751_ ), .Z(\mreg/_06622_ ) );
BUF_X1 \mreg/_13612_ ( .A(\mreg/_00752_ ), .Z(\mreg/_06623_ ) );
BUF_X1 \mreg/_13613_ ( .A(\mreg/_00753_ ), .Z(\mreg/_06624_ ) );
BUF_X1 \mreg/_13614_ ( .A(\mreg/_00754_ ), .Z(\mreg/_06625_ ) );
BUF_X1 \mreg/_13615_ ( .A(\mreg/_00755_ ), .Z(\mreg/_06626_ ) );
BUF_X1 \mreg/_13616_ ( .A(\mreg/_00756_ ), .Z(\mreg/_06627_ ) );
BUF_X1 \mreg/_13617_ ( .A(\mreg/_00757_ ), .Z(\mreg/_06628_ ) );
BUF_X1 \mreg/_13618_ ( .A(\mreg/_00758_ ), .Z(\mreg/_06629_ ) );
BUF_X1 \mreg/_13619_ ( .A(\mreg/_00759_ ), .Z(\mreg/_06630_ ) );
BUF_X1 \mreg/_13620_ ( .A(\mreg/_00760_ ), .Z(\mreg/_06631_ ) );
BUF_X1 \mreg/_13621_ ( .A(\mreg/_00761_ ), .Z(\mreg/_06632_ ) );
BUF_X1 \mreg/_13622_ ( .A(\mreg/_00762_ ), .Z(\mreg/_06633_ ) );
BUF_X1 \mreg/_13623_ ( .A(\mreg/_00763_ ), .Z(\mreg/_06634_ ) );
BUF_X1 \mreg/_13624_ ( .A(\mreg/_00764_ ), .Z(\mreg/_06635_ ) );
BUF_X1 \mreg/_13625_ ( .A(\mreg/_00765_ ), .Z(\mreg/_06636_ ) );
BUF_X1 \mreg/_13626_ ( .A(\mreg/_00766_ ), .Z(\mreg/_06637_ ) );
BUF_X1 \mreg/_13627_ ( .A(\mreg/_00767_ ), .Z(\mreg/_06638_ ) );
BUF_X1 \mreg/_13628_ ( .A(\mreg/_00768_ ), .Z(\mreg/_06639_ ) );
BUF_X1 \mreg/_13629_ ( .A(\mreg/_00769_ ), .Z(\mreg/_06640_ ) );
BUF_X1 \mreg/_13630_ ( .A(\mreg/_00770_ ), .Z(\mreg/_06641_ ) );
BUF_X1 \mreg/_13631_ ( .A(\mreg/_00771_ ), .Z(\mreg/_06642_ ) );
BUF_X1 \mreg/_13632_ ( .A(\mreg/_00772_ ), .Z(\mreg/_06643_ ) );
BUF_X1 \mreg/_13633_ ( .A(\mreg/_00773_ ), .Z(\mreg/_06644_ ) );
BUF_X1 \mreg/_13634_ ( .A(\mreg/_00774_ ), .Z(\mreg/_06645_ ) );
BUF_X1 \mreg/_13635_ ( .A(\mreg/_00775_ ), .Z(\mreg/_06646_ ) );
BUF_X1 \mreg/_13636_ ( .A(\mreg/_00776_ ), .Z(\mreg/_06647_ ) );
BUF_X1 \mreg/_13637_ ( .A(\mreg/_00777_ ), .Z(\mreg/_06648_ ) );
BUF_X1 \mreg/_13638_ ( .A(\mreg/_00778_ ), .Z(\mreg/_06649_ ) );
BUF_X1 \mreg/_13639_ ( .A(\mreg/_00779_ ), .Z(\mreg/_06650_ ) );
BUF_X1 \mreg/_13640_ ( .A(\mreg/_00780_ ), .Z(\mreg/_06651_ ) );
BUF_X1 \mreg/_13641_ ( .A(\mreg/_00781_ ), .Z(\mreg/_06652_ ) );
BUF_X1 \mreg/_13642_ ( .A(\mreg/_00782_ ), .Z(\mreg/_06653_ ) );
BUF_X1 \mreg/_13643_ ( .A(\mreg/_00783_ ), .Z(\mreg/_06654_ ) );
BUF_X1 \mreg/_13644_ ( .A(\mreg/_00784_ ), .Z(\mreg/_06655_ ) );
BUF_X1 \mreg/_13645_ ( .A(\mreg/_00785_ ), .Z(\mreg/_06656_ ) );
BUF_X1 \mreg/_13646_ ( .A(\mreg/_00786_ ), .Z(\mreg/_06657_ ) );
BUF_X1 \mreg/_13647_ ( .A(\mreg/_00787_ ), .Z(\mreg/_06658_ ) );
BUF_X1 \mreg/_13648_ ( .A(\mreg/_00788_ ), .Z(\mreg/_06659_ ) );
BUF_X1 \mreg/_13649_ ( .A(\mreg/_00789_ ), .Z(\mreg/_06660_ ) );
BUF_X1 \mreg/_13650_ ( .A(\mreg/_00790_ ), .Z(\mreg/_06661_ ) );
BUF_X1 \mreg/_13651_ ( .A(\mreg/_00791_ ), .Z(\mreg/_06662_ ) );
BUF_X1 \mreg/_13652_ ( .A(\mreg/_00792_ ), .Z(\mreg/_06663_ ) );
BUF_X1 \mreg/_13653_ ( .A(\mreg/_00793_ ), .Z(\mreg/_06664_ ) );
BUF_X1 \mreg/_13654_ ( .A(\mreg/_00794_ ), .Z(\mreg/_06665_ ) );
BUF_X1 \mreg/_13655_ ( .A(\mreg/_00795_ ), .Z(\mreg/_06666_ ) );
BUF_X1 \mreg/_13656_ ( .A(\mreg/_00796_ ), .Z(\mreg/_06667_ ) );
BUF_X1 \mreg/_13657_ ( .A(\mreg/_00797_ ), .Z(\mreg/_06668_ ) );
BUF_X1 \mreg/_13658_ ( .A(\mreg/_00798_ ), .Z(\mreg/_06669_ ) );
BUF_X1 \mreg/_13659_ ( .A(\mreg/_00799_ ), .Z(\mreg/_06670_ ) );
BUF_X1 \mreg/_13660_ ( .A(\mreg/_00800_ ), .Z(\mreg/_06671_ ) );
BUF_X1 \mreg/_13661_ ( .A(\mreg/_00801_ ), .Z(\mreg/_06672_ ) );
BUF_X1 \mreg/_13662_ ( .A(\mreg/_00802_ ), .Z(\mreg/_06673_ ) );
BUF_X1 \mreg/_13663_ ( .A(\mreg/_00803_ ), .Z(\mreg/_06674_ ) );
BUF_X1 \mreg/_13664_ ( .A(\mreg/_00804_ ), .Z(\mreg/_06675_ ) );
BUF_X1 \mreg/_13665_ ( .A(\mreg/_00805_ ), .Z(\mreg/_06676_ ) );
BUF_X1 \mreg/_13666_ ( .A(\mreg/_00806_ ), .Z(\mreg/_06677_ ) );
BUF_X1 \mreg/_13667_ ( .A(\mreg/_00807_ ), .Z(\mreg/_06678_ ) );
BUF_X1 \mreg/_13668_ ( .A(\mreg/_00808_ ), .Z(\mreg/_06679_ ) );
BUF_X1 \mreg/_13669_ ( .A(\mreg/_00809_ ), .Z(\mreg/_06680_ ) );
BUF_X1 \mreg/_13670_ ( .A(\mreg/_00810_ ), .Z(\mreg/_06681_ ) );
BUF_X1 \mreg/_13671_ ( .A(\mreg/_00811_ ), .Z(\mreg/_06682_ ) );
BUF_X1 \mreg/_13672_ ( .A(\mreg/_00812_ ), .Z(\mreg/_06683_ ) );
BUF_X1 \mreg/_13673_ ( .A(\mreg/_00813_ ), .Z(\mreg/_06684_ ) );
BUF_X1 \mreg/_13674_ ( .A(\mreg/_00814_ ), .Z(\mreg/_06685_ ) );
BUF_X1 \mreg/_13675_ ( .A(\mreg/_00815_ ), .Z(\mreg/_06686_ ) );
BUF_X1 \mreg/_13676_ ( .A(\mreg/_00816_ ), .Z(\mreg/_06687_ ) );
BUF_X1 \mreg/_13677_ ( .A(\mreg/_00817_ ), .Z(\mreg/_06688_ ) );
BUF_X1 \mreg/_13678_ ( .A(\mreg/_00818_ ), .Z(\mreg/_06689_ ) );
BUF_X1 \mreg/_13679_ ( .A(\mreg/_00819_ ), .Z(\mreg/_06690_ ) );
BUF_X1 \mreg/_13680_ ( .A(\mreg/_00820_ ), .Z(\mreg/_06691_ ) );
BUF_X1 \mreg/_13681_ ( .A(\mreg/_00821_ ), .Z(\mreg/_06692_ ) );
BUF_X1 \mreg/_13682_ ( .A(\mreg/_00822_ ), .Z(\mreg/_06693_ ) );
BUF_X1 \mreg/_13683_ ( .A(\mreg/_00823_ ), .Z(\mreg/_06694_ ) );
BUF_X1 \mreg/_13684_ ( .A(\mreg/_00824_ ), .Z(\mreg/_06695_ ) );
BUF_X1 \mreg/_13685_ ( .A(\mreg/_00825_ ), .Z(\mreg/_06696_ ) );
BUF_X1 \mreg/_13686_ ( .A(\mreg/_00826_ ), .Z(\mreg/_06697_ ) );
BUF_X1 \mreg/_13687_ ( .A(\mreg/_00827_ ), .Z(\mreg/_06698_ ) );
BUF_X1 \mreg/_13688_ ( .A(\mreg/_00828_ ), .Z(\mreg/_06699_ ) );
BUF_X1 \mreg/_13689_ ( .A(\mreg/_00829_ ), .Z(\mreg/_06700_ ) );
BUF_X1 \mreg/_13690_ ( .A(\mreg/_00830_ ), .Z(\mreg/_06701_ ) );
BUF_X1 \mreg/_13691_ ( .A(\mreg/_00831_ ), .Z(\mreg/_06702_ ) );
BUF_X1 \mreg/_13692_ ( .A(\mreg/_00832_ ), .Z(\mreg/_06703_ ) );
BUF_X1 \mreg/_13693_ ( .A(\mreg/_00833_ ), .Z(\mreg/_06704_ ) );
BUF_X1 \mreg/_13694_ ( .A(\mreg/_00834_ ), .Z(\mreg/_06705_ ) );
BUF_X1 \mreg/_13695_ ( .A(\mreg/_00835_ ), .Z(\mreg/_06706_ ) );
BUF_X1 \mreg/_13696_ ( .A(\mreg/_00836_ ), .Z(\mreg/_06707_ ) );
BUF_X1 \mreg/_13697_ ( .A(\mreg/_00837_ ), .Z(\mreg/_06708_ ) );
BUF_X1 \mreg/_13698_ ( .A(\mreg/_00838_ ), .Z(\mreg/_06709_ ) );
BUF_X1 \mreg/_13699_ ( .A(\mreg/_00839_ ), .Z(\mreg/_06710_ ) );
BUF_X1 \mreg/_13700_ ( .A(\mreg/_00840_ ), .Z(\mreg/_06711_ ) );
BUF_X1 \mreg/_13701_ ( .A(\mreg/_00841_ ), .Z(\mreg/_06712_ ) );
BUF_X1 \mreg/_13702_ ( .A(\mreg/_00842_ ), .Z(\mreg/_06713_ ) );
BUF_X1 \mreg/_13703_ ( .A(\mreg/_00843_ ), .Z(\mreg/_06714_ ) );
BUF_X1 \mreg/_13704_ ( .A(\mreg/_00844_ ), .Z(\mreg/_06715_ ) );
BUF_X1 \mreg/_13705_ ( .A(\mreg/_00845_ ), .Z(\mreg/_06716_ ) );
BUF_X1 \mreg/_13706_ ( .A(\mreg/_00846_ ), .Z(\mreg/_06717_ ) );
BUF_X1 \mreg/_13707_ ( .A(\mreg/_00847_ ), .Z(\mreg/_06718_ ) );
BUF_X1 \mreg/_13708_ ( .A(\mreg/_00848_ ), .Z(\mreg/_06719_ ) );
BUF_X1 \mreg/_13709_ ( .A(\mreg/_00849_ ), .Z(\mreg/_06720_ ) );
BUF_X1 \mreg/_13710_ ( .A(\mreg/_00850_ ), .Z(\mreg/_06721_ ) );
BUF_X1 \mreg/_13711_ ( .A(\mreg/_00851_ ), .Z(\mreg/_06722_ ) );
BUF_X1 \mreg/_13712_ ( .A(\mreg/_00852_ ), .Z(\mreg/_06723_ ) );
BUF_X1 \mreg/_13713_ ( .A(\mreg/_00853_ ), .Z(\mreg/_06724_ ) );
BUF_X1 \mreg/_13714_ ( .A(\mreg/_00854_ ), .Z(\mreg/_06725_ ) );
BUF_X1 \mreg/_13715_ ( .A(\mreg/_00855_ ), .Z(\mreg/_06726_ ) );
BUF_X1 \mreg/_13716_ ( .A(\mreg/_00856_ ), .Z(\mreg/_06727_ ) );
BUF_X1 \mreg/_13717_ ( .A(\mreg/_00857_ ), .Z(\mreg/_06728_ ) );
BUF_X1 \mreg/_13718_ ( .A(\mreg/_00858_ ), .Z(\mreg/_06729_ ) );
BUF_X1 \mreg/_13719_ ( .A(\mreg/_00859_ ), .Z(\mreg/_06730_ ) );
BUF_X1 \mreg/_13720_ ( .A(\mreg/_00860_ ), .Z(\mreg/_06731_ ) );
BUF_X1 \mreg/_13721_ ( .A(\mreg/_00861_ ), .Z(\mreg/_06732_ ) );
BUF_X1 \mreg/_13722_ ( .A(\mreg/_00862_ ), .Z(\mreg/_06733_ ) );
BUF_X1 \mreg/_13723_ ( .A(\mreg/_00863_ ), .Z(\mreg/_06734_ ) );
BUF_X1 \mreg/_13724_ ( .A(\mreg/_00864_ ), .Z(\mreg/_06735_ ) );
BUF_X1 \mreg/_13725_ ( .A(\mreg/_00865_ ), .Z(\mreg/_06736_ ) );
BUF_X1 \mreg/_13726_ ( .A(\mreg/_00866_ ), .Z(\mreg/_06737_ ) );
BUF_X1 \mreg/_13727_ ( .A(\mreg/_00867_ ), .Z(\mreg/_06738_ ) );
BUF_X1 \mreg/_13728_ ( .A(\mreg/_00868_ ), .Z(\mreg/_06739_ ) );
BUF_X1 \mreg/_13729_ ( .A(\mreg/_00869_ ), .Z(\mreg/_06740_ ) );
BUF_X1 \mreg/_13730_ ( .A(\mreg/_00870_ ), .Z(\mreg/_06741_ ) );
BUF_X1 \mreg/_13731_ ( .A(\mreg/_00871_ ), .Z(\mreg/_06742_ ) );
BUF_X1 \mreg/_13732_ ( .A(\mreg/_00872_ ), .Z(\mreg/_06743_ ) );
BUF_X1 \mreg/_13733_ ( .A(\mreg/_00873_ ), .Z(\mreg/_06744_ ) );
BUF_X1 \mreg/_13734_ ( .A(\mreg/_00874_ ), .Z(\mreg/_06745_ ) );
BUF_X1 \mreg/_13735_ ( .A(\mreg/_00875_ ), .Z(\mreg/_06746_ ) );
BUF_X1 \mreg/_13736_ ( .A(\mreg/_00876_ ), .Z(\mreg/_06747_ ) );
BUF_X1 \mreg/_13737_ ( .A(\mreg/_00877_ ), .Z(\mreg/_06748_ ) );
BUF_X1 \mreg/_13738_ ( .A(\mreg/_00878_ ), .Z(\mreg/_06749_ ) );
BUF_X1 \mreg/_13739_ ( .A(\mreg/_00879_ ), .Z(\mreg/_06750_ ) );
BUF_X1 \mreg/_13740_ ( .A(\mreg/_00880_ ), .Z(\mreg/_06751_ ) );
BUF_X1 \mreg/_13741_ ( .A(\mreg/_00881_ ), .Z(\mreg/_06752_ ) );
BUF_X1 \mreg/_13742_ ( .A(\mreg/_00882_ ), .Z(\mreg/_06753_ ) );
BUF_X1 \mreg/_13743_ ( .A(\mreg/_00883_ ), .Z(\mreg/_06754_ ) );
BUF_X1 \mreg/_13744_ ( .A(\mreg/_00884_ ), .Z(\mreg/_06755_ ) );
BUF_X1 \mreg/_13745_ ( .A(\mreg/_00885_ ), .Z(\mreg/_06756_ ) );
BUF_X1 \mreg/_13746_ ( .A(\mreg/_00886_ ), .Z(\mreg/_06757_ ) );
BUF_X1 \mreg/_13747_ ( .A(\mreg/_00887_ ), .Z(\mreg/_06758_ ) );
BUF_X1 \mreg/_13748_ ( .A(\mreg/_00888_ ), .Z(\mreg/_06759_ ) );
BUF_X1 \mreg/_13749_ ( .A(\mreg/_00889_ ), .Z(\mreg/_06760_ ) );
BUF_X1 \mreg/_13750_ ( .A(\mreg/_00890_ ), .Z(\mreg/_06761_ ) );
BUF_X1 \mreg/_13751_ ( .A(\mreg/_00891_ ), .Z(\mreg/_06762_ ) );
BUF_X1 \mreg/_13752_ ( .A(\mreg/_00892_ ), .Z(\mreg/_06763_ ) );
BUF_X1 \mreg/_13753_ ( .A(\mreg/_00893_ ), .Z(\mreg/_06764_ ) );
BUF_X1 \mreg/_13754_ ( .A(\mreg/_00894_ ), .Z(\mreg/_06765_ ) );
BUF_X1 \mreg/_13755_ ( .A(\mreg/_00895_ ), .Z(\mreg/_06766_ ) );
BUF_X1 \mreg/_13756_ ( .A(\mreg/_00896_ ), .Z(\mreg/_06767_ ) );
BUF_X1 \mreg/_13757_ ( .A(\mreg/_00897_ ), .Z(\mreg/_06768_ ) );
BUF_X1 \mreg/_13758_ ( .A(\mreg/_00898_ ), .Z(\mreg/_06769_ ) );
BUF_X1 \mreg/_13759_ ( .A(\mreg/_00899_ ), .Z(\mreg/_06770_ ) );
BUF_X1 \mreg/_13760_ ( .A(\mreg/_00900_ ), .Z(\mreg/_06771_ ) );
BUF_X1 \mreg/_13761_ ( .A(\mreg/_00901_ ), .Z(\mreg/_06772_ ) );
BUF_X1 \mreg/_13762_ ( .A(\mreg/_00902_ ), .Z(\mreg/_06773_ ) );
BUF_X1 \mreg/_13763_ ( .A(\mreg/_00903_ ), .Z(\mreg/_06774_ ) );
BUF_X1 \mreg/_13764_ ( .A(\mreg/_00904_ ), .Z(\mreg/_06775_ ) );
BUF_X1 \mreg/_13765_ ( .A(\mreg/_00905_ ), .Z(\mreg/_06776_ ) );
BUF_X1 \mreg/_13766_ ( .A(\mreg/_00906_ ), .Z(\mreg/_06777_ ) );
BUF_X1 \mreg/_13767_ ( .A(\mreg/_00907_ ), .Z(\mreg/_06778_ ) );
BUF_X1 \mreg/_13768_ ( .A(\mreg/_00908_ ), .Z(\mreg/_06779_ ) );
BUF_X1 \mreg/_13769_ ( .A(\mreg/_00909_ ), .Z(\mreg/_06780_ ) );
BUF_X1 \mreg/_13770_ ( .A(\mreg/_00910_ ), .Z(\mreg/_06781_ ) );
BUF_X1 \mreg/_13771_ ( .A(\mreg/_00911_ ), .Z(\mreg/_06782_ ) );
BUF_X1 \mreg/_13772_ ( .A(\mreg/_00912_ ), .Z(\mreg/_06783_ ) );
BUF_X1 \mreg/_13773_ ( .A(\mreg/_00913_ ), .Z(\mreg/_06784_ ) );
BUF_X1 \mreg/_13774_ ( .A(\mreg/_00914_ ), .Z(\mreg/_06785_ ) );
BUF_X1 \mreg/_13775_ ( .A(\mreg/_00915_ ), .Z(\mreg/_06786_ ) );
BUF_X1 \mreg/_13776_ ( .A(\mreg/_00916_ ), .Z(\mreg/_06787_ ) );
BUF_X1 \mreg/_13777_ ( .A(\mreg/_00917_ ), .Z(\mreg/_06788_ ) );
BUF_X1 \mreg/_13778_ ( .A(\mreg/_00918_ ), .Z(\mreg/_06789_ ) );
BUF_X1 \mreg/_13779_ ( .A(\mreg/_00919_ ), .Z(\mreg/_06790_ ) );
BUF_X1 \mreg/_13780_ ( .A(\mreg/_00920_ ), .Z(\mreg/_06791_ ) );
BUF_X1 \mreg/_13781_ ( .A(\mreg/_00921_ ), .Z(\mreg/_06792_ ) );
BUF_X1 \mreg/_13782_ ( .A(\mreg/_00922_ ), .Z(\mreg/_06793_ ) );
BUF_X1 \mreg/_13783_ ( .A(\mreg/_00923_ ), .Z(\mreg/_06794_ ) );
BUF_X1 \mreg/_13784_ ( .A(\mreg/_00924_ ), .Z(\mreg/_06795_ ) );
BUF_X1 \mreg/_13785_ ( .A(\mreg/_00925_ ), .Z(\mreg/_06796_ ) );
BUF_X1 \mreg/_13786_ ( .A(\mreg/_00926_ ), .Z(\mreg/_06797_ ) );
BUF_X1 \mreg/_13787_ ( .A(\mreg/_00927_ ), .Z(\mreg/_06798_ ) );
BUF_X1 \mreg/_13788_ ( .A(\mreg/_00928_ ), .Z(\mreg/_06799_ ) );
BUF_X1 \mreg/_13789_ ( .A(\mreg/_00929_ ), .Z(\mreg/_06800_ ) );
BUF_X1 \mreg/_13790_ ( .A(\mreg/_00930_ ), .Z(\mreg/_06801_ ) );
BUF_X1 \mreg/_13791_ ( .A(\mreg/_00931_ ), .Z(\mreg/_06802_ ) );
BUF_X1 \mreg/_13792_ ( .A(\mreg/_00932_ ), .Z(\mreg/_06803_ ) );
BUF_X1 \mreg/_13793_ ( .A(\mreg/_00933_ ), .Z(\mreg/_06804_ ) );
BUF_X1 \mreg/_13794_ ( .A(\mreg/_00934_ ), .Z(\mreg/_06805_ ) );
BUF_X1 \mreg/_13795_ ( .A(\mreg/_00935_ ), .Z(\mreg/_06806_ ) );
BUF_X1 \mreg/_13796_ ( .A(\mreg/_00936_ ), .Z(\mreg/_06807_ ) );
BUF_X1 \mreg/_13797_ ( .A(\mreg/_00937_ ), .Z(\mreg/_06808_ ) );
BUF_X1 \mreg/_13798_ ( .A(\mreg/_00938_ ), .Z(\mreg/_06809_ ) );
BUF_X1 \mreg/_13799_ ( .A(\mreg/_00939_ ), .Z(\mreg/_06810_ ) );
BUF_X1 \mreg/_13800_ ( .A(\mreg/_00940_ ), .Z(\mreg/_06811_ ) );
BUF_X1 \mreg/_13801_ ( .A(\mreg/_00941_ ), .Z(\mreg/_06812_ ) );
BUF_X1 \mreg/_13802_ ( .A(\mreg/_00942_ ), .Z(\mreg/_06813_ ) );
BUF_X1 \mreg/_13803_ ( .A(\mreg/_00943_ ), .Z(\mreg/_06814_ ) );
BUF_X1 \mreg/_13804_ ( .A(\mreg/_00944_ ), .Z(\mreg/_06815_ ) );
BUF_X1 \mreg/_13805_ ( .A(\mreg/_00945_ ), .Z(\mreg/_06816_ ) );
BUF_X1 \mreg/_13806_ ( .A(\mreg/_00946_ ), .Z(\mreg/_06817_ ) );
BUF_X1 \mreg/_13807_ ( .A(\mreg/_00947_ ), .Z(\mreg/_06818_ ) );
BUF_X1 \mreg/_13808_ ( .A(\mreg/_00948_ ), .Z(\mreg/_06819_ ) );
BUF_X1 \mreg/_13809_ ( .A(\mreg/_00949_ ), .Z(\mreg/_06820_ ) );
BUF_X1 \mreg/_13810_ ( .A(\mreg/_00950_ ), .Z(\mreg/_06821_ ) );
BUF_X1 \mreg/_13811_ ( .A(\mreg/_00951_ ), .Z(\mreg/_06822_ ) );
BUF_X1 \mreg/_13812_ ( .A(\mreg/_00952_ ), .Z(\mreg/_06823_ ) );
BUF_X1 \mreg/_13813_ ( .A(\mreg/_00953_ ), .Z(\mreg/_06824_ ) );
BUF_X1 \mreg/_13814_ ( .A(\mreg/_00954_ ), .Z(\mreg/_06825_ ) );
BUF_X1 \mreg/_13815_ ( .A(\mreg/_00955_ ), .Z(\mreg/_06826_ ) );
BUF_X1 \mreg/_13816_ ( .A(\mreg/_00956_ ), .Z(\mreg/_06827_ ) );
BUF_X1 \mreg/_13817_ ( .A(\mreg/_00957_ ), .Z(\mreg/_06828_ ) );
BUF_X1 \mreg/_13818_ ( .A(\mreg/_00958_ ), .Z(\mreg/_06829_ ) );
BUF_X1 \mreg/_13819_ ( .A(\mreg/_00959_ ), .Z(\mreg/_06830_ ) );
BUF_X1 \mreg/_13820_ ( .A(\mreg/_00960_ ), .Z(\mreg/_06831_ ) );
BUF_X1 \mreg/_13821_ ( .A(\mreg/_00961_ ), .Z(\mreg/_06832_ ) );
BUF_X1 \mreg/_13822_ ( .A(\mreg/_00962_ ), .Z(\mreg/_06833_ ) );
BUF_X1 \mreg/_13823_ ( .A(\mreg/_00963_ ), .Z(\mreg/_06834_ ) );
BUF_X1 \mreg/_13824_ ( .A(\mreg/_00964_ ), .Z(\mreg/_06835_ ) );
BUF_X1 \mreg/_13825_ ( .A(\mreg/_00965_ ), .Z(\mreg/_06836_ ) );
BUF_X1 \mreg/_13826_ ( .A(\mreg/_00966_ ), .Z(\mreg/_06837_ ) );
BUF_X1 \mreg/_13827_ ( .A(\mreg/_00967_ ), .Z(\mreg/_06838_ ) );
BUF_X1 \mreg/_13828_ ( .A(\mreg/_00968_ ), .Z(\mreg/_06839_ ) );
BUF_X1 \mreg/_13829_ ( .A(\mreg/_00969_ ), .Z(\mreg/_06840_ ) );
BUF_X1 \mreg/_13830_ ( .A(\mreg/_00970_ ), .Z(\mreg/_06841_ ) );
BUF_X1 \mreg/_13831_ ( .A(\mreg/_00971_ ), .Z(\mreg/_06842_ ) );
BUF_X1 \mreg/_13832_ ( .A(\mreg/_00972_ ), .Z(\mreg/_06843_ ) );
BUF_X1 \mreg/_13833_ ( .A(\mreg/_00973_ ), .Z(\mreg/_06844_ ) );
BUF_X1 \mreg/_13834_ ( .A(\mreg/_00974_ ), .Z(\mreg/_06845_ ) );
BUF_X1 \mreg/_13835_ ( .A(\mreg/_00975_ ), .Z(\mreg/_06846_ ) );
BUF_X1 \mreg/_13836_ ( .A(\mreg/_00976_ ), .Z(\mreg/_06847_ ) );
BUF_X1 \mreg/_13837_ ( .A(\mreg/_00977_ ), .Z(\mreg/_06848_ ) );
BUF_X1 \mreg/_13838_ ( .A(\mreg/_00978_ ), .Z(\mreg/_06849_ ) );
BUF_X1 \mreg/_13839_ ( .A(\mreg/_00979_ ), .Z(\mreg/_06850_ ) );
BUF_X1 \mreg/_13840_ ( .A(\mreg/_00980_ ), .Z(\mreg/_06851_ ) );
BUF_X1 \mreg/_13841_ ( .A(\mreg/_00981_ ), .Z(\mreg/_06852_ ) );
BUF_X1 \mreg/_13842_ ( .A(\mreg/_00982_ ), .Z(\mreg/_06853_ ) );
BUF_X1 \mreg/_13843_ ( .A(\mreg/_00983_ ), .Z(\mreg/_06854_ ) );
BUF_X1 \mreg/_13844_ ( .A(\mreg/_00984_ ), .Z(\mreg/_06855_ ) );
BUF_X1 \mreg/_13845_ ( .A(\mreg/_00985_ ), .Z(\mreg/_06856_ ) );
BUF_X1 \mreg/_13846_ ( .A(\mreg/_00986_ ), .Z(\mreg/_06857_ ) );
BUF_X1 \mreg/_13847_ ( .A(\mreg/_00987_ ), .Z(\mreg/_06858_ ) );
BUF_X1 \mreg/_13848_ ( .A(\mreg/_00988_ ), .Z(\mreg/_06859_ ) );
BUF_X1 \mreg/_13849_ ( .A(\mreg/_00989_ ), .Z(\mreg/_06860_ ) );
BUF_X1 \mreg/_13850_ ( .A(\mreg/_00990_ ), .Z(\mreg/_06861_ ) );
BUF_X1 \mreg/_13851_ ( .A(\mreg/_00991_ ), .Z(\mreg/_06862_ ) );
BUF_X1 \mreg/_13852_ ( .A(\mreg/_00992_ ), .Z(\mreg/_06863_ ) );
BUF_X1 \mreg/_13853_ ( .A(\mreg/_00993_ ), .Z(\mreg/_06864_ ) );
BUF_X1 \mreg/_13854_ ( .A(\mreg/_00994_ ), .Z(\mreg/_06865_ ) );
BUF_X1 \mreg/_13855_ ( .A(\mreg/_00995_ ), .Z(\mreg/_06866_ ) );
BUF_X1 \mreg/_13856_ ( .A(\mreg/_00996_ ), .Z(\mreg/_06867_ ) );
BUF_X1 \mreg/_13857_ ( .A(\mreg/_00997_ ), .Z(\mreg/_06868_ ) );
BUF_X1 \mreg/_13858_ ( .A(\mreg/_00998_ ), .Z(\mreg/_06869_ ) );
BUF_X1 \mreg/_13859_ ( .A(\mreg/_00999_ ), .Z(\mreg/_06870_ ) );
BUF_X1 \mreg/_13860_ ( .A(\mreg/_01000_ ), .Z(\mreg/_06871_ ) );
BUF_X1 \mreg/_13861_ ( .A(\mreg/_01001_ ), .Z(\mreg/_06872_ ) );
BUF_X1 \mreg/_13862_ ( .A(\mreg/_01002_ ), .Z(\mreg/_06873_ ) );
BUF_X1 \mreg/_13863_ ( .A(\mreg/_01003_ ), .Z(\mreg/_06874_ ) );
BUF_X1 \mreg/_13864_ ( .A(\mreg/_01004_ ), .Z(\mreg/_06875_ ) );
BUF_X1 \mreg/_13865_ ( .A(\mreg/_01005_ ), .Z(\mreg/_06876_ ) );
BUF_X1 \mreg/_13866_ ( .A(\mreg/_01006_ ), .Z(\mreg/_06877_ ) );
BUF_X1 \mreg/_13867_ ( .A(\mreg/_01007_ ), .Z(\mreg/_06878_ ) );
BUF_X1 \mreg/_13868_ ( .A(\mreg/_01008_ ), .Z(\mreg/_06879_ ) );
BUF_X1 \mreg/_13869_ ( .A(\mreg/_01009_ ), .Z(\mreg/_06880_ ) );
BUF_X1 \mreg/_13870_ ( .A(\mreg/_01010_ ), .Z(\mreg/_06881_ ) );
BUF_X1 \mreg/_13871_ ( .A(\mreg/_01011_ ), .Z(\mreg/_06882_ ) );
BUF_X1 \mreg/_13872_ ( .A(\mreg/_01012_ ), .Z(\mreg/_06883_ ) );
BUF_X1 \mreg/_13873_ ( .A(\mreg/_01013_ ), .Z(\mreg/_06884_ ) );
BUF_X1 \mreg/_13874_ ( .A(\mreg/_01014_ ), .Z(\mreg/_06885_ ) );
BUF_X1 \mreg/_13875_ ( .A(\mreg/_01015_ ), .Z(\mreg/_06886_ ) );
BUF_X1 \mreg/_13876_ ( .A(\mreg/_01016_ ), .Z(\mreg/_06887_ ) );
BUF_X1 \mreg/_13877_ ( .A(\mreg/_01017_ ), .Z(\mreg/_06888_ ) );
BUF_X1 \mreg/_13878_ ( .A(\mreg/_01018_ ), .Z(\mreg/_06889_ ) );
BUF_X1 \mreg/_13879_ ( .A(\mreg/_01019_ ), .Z(\mreg/_06890_ ) );
BUF_X1 \mreg/_13880_ ( .A(\mreg/_01020_ ), .Z(\mreg/_06891_ ) );
BUF_X1 \mreg/_13881_ ( .A(\mreg/_01021_ ), .Z(\mreg/_06892_ ) );
BUF_X1 \mreg/_13882_ ( .A(\mreg/_01022_ ), .Z(\mreg/_06893_ ) );
BUF_X1 \mreg/_13883_ ( .A(\mreg/_01023_ ), .Z(\mreg/_06894_ ) );
BUF_X1 \mreg/_13884_ ( .A(\mreg/_01024_ ), .Z(\mreg/_06895_ ) );
BUF_X1 \mreg/_13885_ ( .A(\mreg/_01025_ ), .Z(\mreg/_06896_ ) );
BUF_X1 \mreg/_13886_ ( .A(\mreg/_01026_ ), .Z(\mreg/_06897_ ) );
BUF_X1 \mreg/_13887_ ( .A(\mreg/_01027_ ), .Z(\mreg/_06898_ ) );
BUF_X1 \mreg/_13888_ ( .A(\mreg/_01028_ ), .Z(\mreg/_06899_ ) );
BUF_X1 \mreg/_13889_ ( .A(\mreg/_01029_ ), .Z(\mreg/_06900_ ) );
BUF_X1 \mreg/_13890_ ( .A(\mreg/_01030_ ), .Z(\mreg/_06901_ ) );
BUF_X1 \mreg/_13891_ ( .A(\mreg/_01031_ ), .Z(\mreg/_06902_ ) );
BUF_X1 \mreg/_13892_ ( .A(\mreg/_01032_ ), .Z(\mreg/_06903_ ) );
BUF_X1 \mreg/_13893_ ( .A(\mreg/_01033_ ), .Z(\mreg/_06904_ ) );
BUF_X1 \mreg/_13894_ ( .A(\mreg/_01034_ ), .Z(\mreg/_06905_ ) );
BUF_X1 \mreg/_13895_ ( .A(\mreg/_01035_ ), .Z(\mreg/_06906_ ) );
BUF_X1 \mreg/_13896_ ( .A(\mreg/_01036_ ), .Z(\mreg/_06907_ ) );
BUF_X1 \mreg/_13897_ ( .A(\mreg/_01037_ ), .Z(\mreg/_06908_ ) );
BUF_X1 \mreg/_13898_ ( .A(\mreg/_01038_ ), .Z(\mreg/_06909_ ) );
BUF_X1 \mreg/_13899_ ( .A(\mreg/_01039_ ), .Z(\mreg/_06910_ ) );
BUF_X1 \mreg/_13900_ ( .A(\mreg/_01040_ ), .Z(\mreg/_06911_ ) );
BUF_X1 \mreg/_13901_ ( .A(\mreg/_01041_ ), .Z(\mreg/_06912_ ) );
BUF_X1 \mreg/_13902_ ( .A(\mreg/_01042_ ), .Z(\mreg/_06913_ ) );
BUF_X1 \mreg/_13903_ ( .A(\mreg/_01043_ ), .Z(\mreg/_06914_ ) );
BUF_X1 \mreg/_13904_ ( .A(\mreg/_01044_ ), .Z(\mreg/_06915_ ) );
BUF_X1 \mreg/_13905_ ( .A(\mreg/_01045_ ), .Z(\mreg/_06916_ ) );
BUF_X1 \mreg/_13906_ ( .A(\mreg/_01046_ ), .Z(\mreg/_06917_ ) );
BUF_X1 \mreg/_13907_ ( .A(\mreg/_01047_ ), .Z(\mreg/_06918_ ) );
BUF_X1 \mreg/_13908_ ( .A(\mreg/_01048_ ), .Z(\mreg/_06919_ ) );
BUF_X1 \mreg/_13909_ ( .A(\mreg/_01049_ ), .Z(\mreg/_06920_ ) );
BUF_X1 \mreg/_13910_ ( .A(\mreg/_01050_ ), .Z(\mreg/_06921_ ) );
BUF_X1 \mreg/_13911_ ( .A(\mreg/_01051_ ), .Z(\mreg/_06922_ ) );
BUF_X1 \mreg/_13912_ ( .A(\mreg/_01052_ ), .Z(\mreg/_06923_ ) );
BUF_X1 \mreg/_13913_ ( .A(\mreg/_01053_ ), .Z(\mreg/_06924_ ) );
INV_X1 \msram/_15_ ( .A(\msram/_01_ ), .ZN(\msram/_07_ ) );
NOR3_X1 \msram/_16_ ( .A1(\msram/_07_ ), .A2(\msram/_00_ ), .A3(\msram/_08_ ), .ZN(\msram/_02_ ) );
NAND2_X1 \msram/_17_ ( .A1(\msram/_05_ ), .A2(\msram/_09_ ), .ZN(\msram/_06_ ) );
NOR3_X1 \msram/_18_ ( .A1(\msram/_06_ ), .A2(\msram/_04_ ), .A3(\msram/_08_ ), .ZN(\msram/_03_ ) );
DFF_X1 \msram/_19_ ( .CK(clk ), .D(\msram/_13_ ), .Q(arready ), .QN(\msram/_11_ ) );
DFF_X1 \msram/_20_ ( .CK(clk ), .D(\msram/_14_ ), .Q(awready ), .QN(\msram/_10_ ) );
LOGIC0_X1 \msram/_21_ ( .Z(\msram/_12_ ) );
BUF_X1 \msram/_22_ ( .A(\msram/_12_ ), .Z(\bresp[0] ) );
BUF_X1 \msram/_23_ ( .A(\msram/_12_ ), .Z(\bresp[1] ) );
BUF_X1 \msram/_24_ ( .A(\msram/_12_ ), .Z(bvalid ) );
BUF_X1 \msram/_25_ ( .A(\msram/_12_ ), .Z(\rdata[0] ) );
BUF_X1 \msram/_26_ ( .A(\msram/_12_ ), .Z(\rdata[1] ) );
BUF_X1 \msram/_27_ ( .A(\msram/_12_ ), .Z(\rdata[2] ) );
BUF_X1 \msram/_28_ ( .A(\msram/_12_ ), .Z(\rdata[3] ) );
BUF_X1 \msram/_29_ ( .A(\msram/_12_ ), .Z(\rdata[4] ) );
BUF_X1 \msram/_30_ ( .A(\msram/_12_ ), .Z(\rdata[5] ) );
BUF_X1 \msram/_31_ ( .A(\msram/_12_ ), .Z(\rdata[6] ) );
BUF_X1 \msram/_32_ ( .A(\msram/_12_ ), .Z(\rdata[7] ) );
BUF_X1 \msram/_33_ ( .A(\msram/_12_ ), .Z(\rdata[8] ) );
BUF_X1 \msram/_34_ ( .A(\msram/_12_ ), .Z(\rdata[9] ) );
BUF_X1 \msram/_35_ ( .A(\msram/_12_ ), .Z(\rdata[10] ) );
BUF_X1 \msram/_36_ ( .A(\msram/_12_ ), .Z(\rdata[11] ) );
BUF_X1 \msram/_37_ ( .A(\msram/_12_ ), .Z(\rdata[12] ) );
BUF_X1 \msram/_38_ ( .A(\msram/_12_ ), .Z(\rdata[13] ) );
BUF_X1 \msram/_39_ ( .A(\msram/_12_ ), .Z(\rdata[14] ) );
BUF_X1 \msram/_40_ ( .A(\msram/_12_ ), .Z(\rdata[15] ) );
BUF_X1 \msram/_41_ ( .A(\msram/_12_ ), .Z(\rdata[16] ) );
BUF_X1 \msram/_42_ ( .A(\msram/_12_ ), .Z(\rdata[17] ) );
BUF_X1 \msram/_43_ ( .A(\msram/_12_ ), .Z(\rdata[18] ) );
BUF_X1 \msram/_44_ ( .A(\msram/_12_ ), .Z(\rdata[19] ) );
BUF_X1 \msram/_45_ ( .A(\msram/_12_ ), .Z(\rdata[20] ) );
BUF_X1 \msram/_46_ ( .A(\msram/_12_ ), .Z(\rdata[21] ) );
BUF_X1 \msram/_47_ ( .A(\msram/_12_ ), .Z(\rdata[22] ) );
BUF_X1 \msram/_48_ ( .A(\msram/_12_ ), .Z(\rdata[23] ) );
BUF_X1 \msram/_49_ ( .A(\msram/_12_ ), .Z(\rdata[24] ) );
BUF_X1 \msram/_50_ ( .A(\msram/_12_ ), .Z(\rdata[25] ) );
BUF_X1 \msram/_51_ ( .A(\msram/_12_ ), .Z(\rdata[26] ) );
BUF_X1 \msram/_52_ ( .A(\msram/_12_ ), .Z(\rdata[27] ) );
BUF_X1 \msram/_53_ ( .A(\msram/_12_ ), .Z(\rdata[28] ) );
BUF_X1 \msram/_54_ ( .A(\msram/_12_ ), .Z(\rdata[29] ) );
BUF_X1 \msram/_55_ ( .A(\msram/_12_ ), .Z(\rdata[30] ) );
BUF_X1 \msram/_56_ ( .A(\msram/_12_ ), .Z(\rdata[31] ) );
BUF_X1 \msram/_57_ ( .A(\msram/_12_ ), .Z(\rresp[0] ) );
BUF_X1 \msram/_58_ ( .A(\msram/_12_ ), .Z(\rresp[1] ) );
BUF_X1 \msram/_59_ ( .A(\msram/_12_ ), .Z(rvalid ) );
BUF_X1 \msram/_60_ ( .A(\msram/_12_ ), .Z(wready ) );
BUF_X1 \msram/_61_ ( .A(arvalid ), .Z(\msram/_01_ ) );
BUF_X1 \msram/_62_ ( .A(arready ), .Z(\msram/_00_ ) );
BUF_X1 \msram/_63_ ( .A(awready ), .Z(\msram/_04_ ) );
BUF_X1 \msram/_64_ ( .A(awvalid ), .Z(\msram/_05_ ) );
BUF_X1 \msram/_65_ ( .A(wvalid ), .Z(\msram/_09_ ) );
BUF_X1 \msram/_66_ ( .A(rst ), .Z(\msram/_08_ ) );
BUF_X1 \msram/_67_ ( .A(\msram/_02_ ), .Z(\msram/_13_ ) );
BUF_X1 \msram/_68_ ( .A(\msram/_03_ ), .Z(\msram/_14_ ) );

endmodule
